module LockingRRArbiter(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [21:0] io_in_0_bits_address,
  input  [31:0] io_in_0_bits_data,
  input  [4:0]  io_in_0_bits_taskID,
  input         io_out_ready,
  output        io_out_valid,
  output [21:0] io_out_bits_address,
  output [31:0] io_out_bits_data,
  output [4:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ,
  output        io_chosen
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? 1'h0 : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_address = io_chosen ? 22'h0 : io_in_0_bits_address; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? 32'h0 : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_out_bits_taskID = io_chosen ? 5'h0 : io_in_0_bits_taskID; // @[Arbiter.scala 42:15]
  assign io_out_bits_Typ = io_chosen ? 8'h0 : 8'h3; // @[Arbiter.scala 42:15]
  assign io_chosen = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 40:13]
endmodule
module ArbiterTree(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [21:0] io_in_0_bits_address,
  input  [31:0] io_in_0_bits_data,
  input  [4:0]  io_in_0_bits_taskID,
  input         io_out_ready,
  output        io_out_valid,
  output [21:0] io_out_bits_address,
  output [31:0] io_out_bits_data,
  output [4:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ
);
  wire  LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_chosen; // @[ArbiterTree.scala 32:13]
  LockingRRArbiter LockingRRArbiter ( // @[ArbiterTree.scala 32:13]
    .io_in_0_ready(LockingRRArbiter_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_io_in_0_valid),
    .io_in_0_bits_address(LockingRRArbiter_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_io_in_0_bits_taskID),
    .io_out_ready(LockingRRArbiter_io_out_ready),
    .io_out_valid(LockingRRArbiter_io_out_valid),
    .io_out_bits_address(LockingRRArbiter_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_io_chosen)
  );
  assign io_in_0_ready = LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_out_valid = LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_address = LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_data = LockingRRArbiter_io_out_bits_data; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_taskID = LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_Typ = LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 65:12]
  assign LockingRRArbiter_io_in_0_valid = io_in_0_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_address = io_in_0_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_data = io_in_0_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_taskID = io_in_0_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_out_ready = io_out_ready; // @[ArbiterTree.scala 65:12]
endmodule
module Arbiter(
  output  io_in_0_ready,
  input   io_in_0_valid,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input   io_out_ready,
  output  io_out_valid
);
  wire  _T; // @[Arbiter.scala 31:78]
  wire  _T_3; // @[Arbiter.scala 135:19]
  assign _T = io_in_0_valid == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_3 = _T == 1'h0; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = _T & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_3 | io_in_1_valid; // @[Arbiter.scala 135:16]
endmodule
module Arbiter_1(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [31:0] io_in_0_bits_data,
  input  [3:0]  io_in_0_bits_mask,
  input  [7:0]  io_in_0_bits_tag,
  input  [4:0]  io_in_0_bits_taskID,
  input         io_in_0_bits_iswrite,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [31:0] io_in_1_bits_data,
  input  [3:0]  io_in_1_bits_mask,
  input  [7:0]  io_in_1_bits_tag,
  input  [4:0]  io_in_1_bits_taskID,
  input         io_in_1_bits_iswrite,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [31:0] io_out_bits_data,
  output [3:0]  io_out_bits_mask,
  output [7:0]  io_out_bits_tag,
  output [4:0]  io_out_bits_taskID,
  output        io_out_bits_iswrite
);
  wire  _T; // @[Arbiter.scala 31:78]
  wire  _T_3; // @[Arbiter.scala 135:19]
  assign _T = io_in_0_valid == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_3 = _T == 1'h0; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = _T & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_3 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_mask = io_in_0_valid ? io_in_0_bits_mask : io_in_1_bits_mask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_tag = io_in_0_valid ? io_in_0_bits_tag : io_in_1_bits_tag; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_taskID = io_in_0_valid ? io_in_0_bits_taskID : io_in_1_bits_taskID; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_iswrite = io_in_0_valid ? io_in_0_bits_iswrite : io_in_1_bits_iswrite; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Demux(
  input         io_en,
  input  [31:0] io_input_data,
  input  [7:0]  io_input_tag,
  input         io_sel,
  output        io_outputs_0_valid,
  output [31:0] io_outputs_0_data,
  output [7:0]  io_outputs_0_tag,
  output        io_outputs_1_valid,
  output [31:0] io_outputs_1_data,
  output [7:0]  io_outputs_1_tag
);
  wire  _GEN_0; // @[Muxes.scala 29:25]
  assign _GEN_0 = 1'h0 == io_sel; // @[Muxes.scala 29:25]
  assign io_outputs_0_valid = io_en & _GEN_0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_0_data = io_input_data; // @[Muxes.scala 23:19]
  assign io_outputs_0_tag = io_input_tag; // @[Muxes.scala 23:19]
  assign io_outputs_1_valid = io_en & io_sel; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_1_data = io_input_data; // @[Muxes.scala 23:19]
  assign io_outputs_1_tag = io_input_tag; // @[Muxes.scala 23:19]
endmodule
module RRArbiter(
  input   clock,
  output  io_in_0_ready,
  input   io_in_0_valid,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input   io_out_ready,
  output  io_out_valid,
  output  io_chosen
);
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Arbiter.scala 67:57]
  wire  _T_5; // @[Arbiter.scala 68:83]
  wire  _T_7; // @[Arbiter.scala 31:68]
  wire  _T_10; // @[Arbiter.scala 31:78]
  wire  _GEN_11; // @[Arbiter.scala 77:27]
  assign _T_3 = 1'h1 > _T_1; // @[Arbiter.scala 67:57]
  assign _T_5 = io_in_1_valid & _T_3; // @[Arbiter.scala 68:83]
  assign _T_7 = _T_5 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_10 = _T_7 == 1'h0; // @[Arbiter.scala 31:78]
  assign _GEN_11 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_5 == 1'h0; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_3 | _T_10; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_chosen = _T_5 | _GEN_11; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_out_valid) begin
      _T_1 <= io_chosen;
    end
  end
endmodule
module Demux_1(
  input   io_en,
  output  io_outputs_0_valid
);
  assign io_outputs_0_valid = io_en; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
endmodule
module DeMuxTree(
  output  io_outputs_0_valid,
  input   io_enable
);
  wire  Demux_io_en; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_0_valid; // @[Muxes.scala 91:13]
  Demux_1 Demux ( // @[Muxes.scala 91:13]
    .io_en(Demux_io_en),
    .io_outputs_0_valid(Demux_io_outputs_0_valid)
  );
  assign io_outputs_0_valid = Demux_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign Demux_io_en = io_enable; // @[Muxes.scala 135:14]
endmodule
module WriteTableEntry(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [21:0] io_NodeReq_bits_address,
  input  [31:0] io_NodeReq_bits_data,
  input  [4:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input         io_output_ready,
  output        io_output_valid,
  output        io_free
);
  reg [4:0] request_R_taskID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_0;
  reg [7:0] sendbytemask; // @[WriteMemoryController.scala 61:29]
  reg [31:0] _RAND_1;
  reg [31:0] ReqAddress; // @[WriteMemoryController.scala 65:27]
  reg [31:0] _RAND_2;
  reg  ptr; // @[WriteMemoryController.scala 70:27]
  reg [31:0] _RAND_3;
  reg [31:0] linebuffer_0; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_4;
  reg [31:0] linebuffer_1; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_5;
  reg [1:0] state; // @[WriteMemoryController.scala 76:68]
  reg [31:0] _RAND_6;
  wire  _T_4; // @[WriteMemoryController.scala 89:21]
  wire [2:0] _T_5; // @[Cat.scala 29:58]
  wire [31:0] _GEN_29; // @[WriteMemoryController.scala 100:37]
  reg  isWrite; // @[WriteMemoryController.scala 108:24]
  reg [31:0] _RAND_7;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire [19:0] _T_10; // @[WriteMemoryController.scala 121:44]
  wire [21:0] _T_11; // @[WriteMemoryController.scala 121:69]
  wire  _T_12; // @[helpers.scala 27:24]
  wire  _T_13; // @[helpers.scala 27:47]
  wire  _T_14; // @[helpers.scala 27:40]
  wire  _T_16; // @[helpers.scala 28:15]
  wire  _T_17; // @[helpers.scala 28:38]
  wire  _T_18; // @[helpers.scala 28:31]
  wire  _T_20; // @[helpers.scala 29:17]
  wire  _T_21; // @[helpers.scala 29:40]
  wire  _T_22; // @[helpers.scala 29:33]
  wire [1:0] _T_28; // @[helpers.scala 39:32]
  wire [4:0] _T_29; // @[Cat.scala 29:58]
  wire [7:0] _T_43; // @[helpers.scala 50:12]
  wire [7:0] _T_44; // @[helpers.scala 49:10]
  wire [7:0] _T_45; // @[helpers.scala 48:19]
  wire [10:0] _GEN_31; // @[helpers.scala 20:26]
  wire [10:0] _T_47; // @[helpers.scala 20:26]
  wire [62:0] _GEN_32; // @[WriteMemoryController.scala 127:41]
  wire [62:0] _T_50; // @[WriteMemoryController.scala 127:41]
  wire [63:0] _T_52;
  wire [31:0] _T_53; // @[WriteMemoryController.scala 127:121]
  wire [31:0] _T_54; // @[WriteMemoryController.scala 127:121]
  wire [10:0] _GEN_10; // @[WriteMemoryController.scala 117:28]
  wire  _T_55; // @[WriteMemoryController.scala 139:15]
  wire  _T_56; // @[WriteMemoryController.scala 139:47]
  wire  _T_57; // @[WriteMemoryController.scala 139:30]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire [3:0] _T_59; // @[WriteMemoryController.scala 144:36]
  wire  _T_61; // @[WriteMemoryController.scala 146:18]
  wire [10:0] _GEN_14; // @[WriteMemoryController.scala 142:29]
  wire [10:0] _GEN_18; // @[WriteMemoryController.scala 139:76]
  wire  _T_62; // @[WriteMemoryController.scala 156:15]
  wire  _T_64; // @[WriteMemoryController.scala 156:32]
  wire  _T_65; // @[WriteMemoryController.scala 158:27]
  wire  _T_68; // @[Decoupled.scala 40:37]
  assign _T_4 = state == 2'h3; // @[WriteMemoryController.scala 89:21]
  assign _T_5 = {ptr,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_29 = {{29'd0}, _T_5}; // @[WriteMemoryController.scala 100:37]
  assign _T_9 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_NodeReq_bits_address[21:2]; // @[WriteMemoryController.scala 121:44]
  assign _T_11 = {_T_10, 2'h0}; // @[WriteMemoryController.scala 121:69]
  assign _T_12 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_13 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_14 = _T_12 | _T_13; // @[helpers.scala 27:40]
  assign _T_16 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_17 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_18 = _T_16 | _T_17; // @[helpers.scala 28:31]
  assign _T_20 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_21 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_22 = _T_20 | _T_21; // @[helpers.scala 29:33]
  assign _T_28 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_29 = {_T_28,3'h0}; // @[Cat.scala 29:58]
  assign _T_43 = _T_22 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_44 = _T_18 ? 8'h1 : _T_43; // @[helpers.scala 49:10]
  assign _T_45 = _T_14 ? 8'h3 : _T_44; // @[helpers.scala 48:19]
  assign _GEN_31 = {{3'd0}, _T_45}; // @[helpers.scala 20:26]
  assign _T_47 = _GEN_31 << _T_28; // @[helpers.scala 20:26]
  assign _GEN_32 = {{31'd0}, io_NodeReq_bits_data}; // @[WriteMemoryController.scala 127:41]
  assign _T_50 = _GEN_32 << _T_29; // @[WriteMemoryController.scala 127:41]
  assign _T_52 = {{1'd0}, _T_50};
  assign _T_53 = _T_52[31:0]; // @[WriteMemoryController.scala 127:121]
  assign _T_54 = _T_52[63:32]; // @[WriteMemoryController.scala 127:121]
  assign _GEN_10 = _T_9 ? _T_47 : {{3'd0}, sendbytemask}; // @[WriteMemoryController.scala 117:28]
  assign _T_55 = state == 2'h1; // @[WriteMemoryController.scala 139:15]
  assign _T_56 = sendbytemask != 8'h0; // @[WriteMemoryController.scala 139:47]
  assign _T_57 = _T_55 & _T_56; // @[WriteMemoryController.scala 139:30]
  assign _T_58 = io_MemReq_ready & io_MemReq_valid; // @[Decoupled.scala 40:37]
  assign _T_59 = sendbytemask[7:4]; // @[WriteMemoryController.scala 144:36]
  assign _T_61 = ptr + 1'h1; // @[WriteMemoryController.scala 146:18]
  assign _GEN_14 = _T_58 ? {{7'd0}, _T_59} : _GEN_10; // @[WriteMemoryController.scala 142:29]
  assign _GEN_18 = _T_57 ? _GEN_14 : _GEN_10; // @[WriteMemoryController.scala 139:76]
  assign _T_62 = state == 2'h2; // @[WriteMemoryController.scala 156:15]
  assign _T_64 = _T_62 & io_MemResp_valid; // @[WriteMemoryController.scala 156:32]
  assign _T_65 = sendbytemask == 8'h0; // @[WriteMemoryController.scala 158:27]
  assign _T_68 = io_output_ready & io_output_valid; // @[Decoupled.scala 40:37]
  assign io_NodeReq_ready = state == 2'h0; // @[WriteMemoryController.scala 87:20]
  assign io_MemReq_valid = _T_55 & _T_56; // @[WriteMemoryController.scala 99:19 WriteMemoryController.scala 140:21]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_29; // @[WriteMemoryController.scala 100:23]
  assign io_MemReq_bits_data = ptr ? linebuffer_1 : linebuffer_0; // @[WriteMemoryController.scala 102:23]
  assign io_MemReq_bits_mask = sendbytemask[3:0]; // @[WriteMemoryController.scala 103:23]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[WriteMemoryController.scala 110:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[WriteMemoryController.scala 109:26]
  assign io_output_valid = state == 2'h3; // @[WriteMemoryController.scala 95:19 WriteMemoryController.scala 168:21]
  assign io_free = state == 2'h0; // @[WriteMemoryController.scala 85:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  request_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  sendbytemask = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ReqAddress = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ptr = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  linebuffer_0 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  linebuffer_1 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  isWrite = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      request_R_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_18[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_9) begin
        ReqAddress <= {{10'd0}, _T_11};
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (_T_4) begin
        ptr <= 1'h0;
      end else begin
        if (_T_57) begin
          if (_T_58) begin
            ptr <= _T_61;
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (_T_9) begin
        linebuffer_0 <= _T_53;
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (_T_9) begin
        linebuffer_1 <= _T_54;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_4) begin
        if (_T_68) begin
          state <= 2'h0;
        end else begin
          if (_T_64) begin
            if (_T_65) begin
              state <= 2'h3;
            end else begin
              state <= 2'h1;
            end
          end else begin
            if (_T_57) begin
              if (_T_58) begin
                state <= 2'h2;
              end else begin
                if (_T_9) begin
                  state <= 2'h1;
                end
              end
            end else begin
              if (_T_9) begin
                state <= 2'h1;
              end
            end
          end
        end
      end else begin
        if (_T_64) begin
          if (_T_65) begin
            state <= 2'h3;
          end else begin
            state <= 2'h1;
          end
        end else begin
          if (_T_57) begin
            if (_T_58) begin
              state <= 2'h2;
            end else begin
              if (_T_9) begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_9) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      isWrite <= 1'h0;
    end else begin
      isWrite <= 1'h1;
    end
  end
endmodule
module WriteTableEntry_1(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [21:0] io_NodeReq_bits_address,
  input  [31:0] io_NodeReq_bits_data,
  input  [4:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input         io_output_ready,
  output        io_output_valid,
  output        io_free
);
  reg  ID; // @[WriteMemoryController.scala 53:32]
  reg [31:0] _RAND_0;
  reg [4:0] request_R_taskID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_1;
  reg [7:0] sendbytemask; // @[WriteMemoryController.scala 61:29]
  reg [31:0] _RAND_2;
  reg [31:0] ReqAddress; // @[WriteMemoryController.scala 65:27]
  reg [31:0] _RAND_3;
  reg  ptr; // @[WriteMemoryController.scala 70:27]
  reg [31:0] _RAND_4;
  reg [31:0] linebuffer_0; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_5;
  reg [31:0] linebuffer_1; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_6;
  reg [1:0] state; // @[WriteMemoryController.scala 76:68]
  reg [31:0] _RAND_7;
  wire  _T_4; // @[WriteMemoryController.scala 89:21]
  wire [2:0] _T_5; // @[Cat.scala 29:58]
  wire [31:0] _GEN_29; // @[WriteMemoryController.scala 100:37]
  reg  myID; // @[WriteMemoryController.scala 106:21]
  reg [31:0] _RAND_8;
  reg  isWrite; // @[WriteMemoryController.scala 108:24]
  reg [31:0] _RAND_9;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire [19:0] _T_10; // @[WriteMemoryController.scala 121:44]
  wire [21:0] _T_11; // @[WriteMemoryController.scala 121:69]
  wire  _T_12; // @[helpers.scala 27:24]
  wire  _T_13; // @[helpers.scala 27:47]
  wire  _T_14; // @[helpers.scala 27:40]
  wire  _T_16; // @[helpers.scala 28:15]
  wire  _T_17; // @[helpers.scala 28:38]
  wire  _T_18; // @[helpers.scala 28:31]
  wire  _T_20; // @[helpers.scala 29:17]
  wire  _T_21; // @[helpers.scala 29:40]
  wire  _T_22; // @[helpers.scala 29:33]
  wire [1:0] _T_28; // @[helpers.scala 39:32]
  wire [4:0] _T_29; // @[Cat.scala 29:58]
  wire [7:0] _T_43; // @[helpers.scala 50:12]
  wire [7:0] _T_44; // @[helpers.scala 49:10]
  wire [7:0] _T_45; // @[helpers.scala 48:19]
  wire [10:0] _GEN_31; // @[helpers.scala 20:26]
  wire [10:0] _T_47; // @[helpers.scala 20:26]
  wire [62:0] _GEN_32; // @[WriteMemoryController.scala 127:41]
  wire [62:0] _T_50; // @[WriteMemoryController.scala 127:41]
  wire [63:0] _T_52;
  wire [31:0] _T_53; // @[WriteMemoryController.scala 127:121]
  wire [31:0] _T_54; // @[WriteMemoryController.scala 127:121]
  wire [10:0] _GEN_10; // @[WriteMemoryController.scala 117:28]
  wire  _T_55; // @[WriteMemoryController.scala 139:15]
  wire  _T_56; // @[WriteMemoryController.scala 139:47]
  wire  _T_57; // @[WriteMemoryController.scala 139:30]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire [3:0] _T_59; // @[WriteMemoryController.scala 144:36]
  wire  _T_61; // @[WriteMemoryController.scala 146:18]
  wire [10:0] _GEN_14; // @[WriteMemoryController.scala 142:29]
  wire [10:0] _GEN_18; // @[WriteMemoryController.scala 139:76]
  wire  _T_62; // @[WriteMemoryController.scala 156:15]
  wire  _T_64; // @[WriteMemoryController.scala 156:32]
  wire  _T_65; // @[WriteMemoryController.scala 158:27]
  wire  _T_68; // @[Decoupled.scala 40:37]
  assign _T_4 = state == 2'h3; // @[WriteMemoryController.scala 89:21]
  assign _T_5 = {ptr,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_29 = {{29'd0}, _T_5}; // @[WriteMemoryController.scala 100:37]
  assign _T_9 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_NodeReq_bits_address[21:2]; // @[WriteMemoryController.scala 121:44]
  assign _T_11 = {_T_10, 2'h0}; // @[WriteMemoryController.scala 121:69]
  assign _T_12 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_13 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_14 = _T_12 | _T_13; // @[helpers.scala 27:40]
  assign _T_16 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_17 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_18 = _T_16 | _T_17; // @[helpers.scala 28:31]
  assign _T_20 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_21 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_22 = _T_20 | _T_21; // @[helpers.scala 29:33]
  assign _T_28 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_29 = {_T_28,3'h0}; // @[Cat.scala 29:58]
  assign _T_43 = _T_22 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_44 = _T_18 ? 8'h1 : _T_43; // @[helpers.scala 49:10]
  assign _T_45 = _T_14 ? 8'h3 : _T_44; // @[helpers.scala 48:19]
  assign _GEN_31 = {{3'd0}, _T_45}; // @[helpers.scala 20:26]
  assign _T_47 = _GEN_31 << _T_28; // @[helpers.scala 20:26]
  assign _GEN_32 = {{31'd0}, io_NodeReq_bits_data}; // @[WriteMemoryController.scala 127:41]
  assign _T_50 = _GEN_32 << _T_29; // @[WriteMemoryController.scala 127:41]
  assign _T_52 = {{1'd0}, _T_50};
  assign _T_53 = _T_52[31:0]; // @[WriteMemoryController.scala 127:121]
  assign _T_54 = _T_52[63:32]; // @[WriteMemoryController.scala 127:121]
  assign _GEN_10 = _T_9 ? _T_47 : {{3'd0}, sendbytemask}; // @[WriteMemoryController.scala 117:28]
  assign _T_55 = state == 2'h1; // @[WriteMemoryController.scala 139:15]
  assign _T_56 = sendbytemask != 8'h0; // @[WriteMemoryController.scala 139:47]
  assign _T_57 = _T_55 & _T_56; // @[WriteMemoryController.scala 139:30]
  assign _T_58 = io_MemReq_ready & io_MemReq_valid; // @[Decoupled.scala 40:37]
  assign _T_59 = sendbytemask[7:4]; // @[WriteMemoryController.scala 144:36]
  assign _T_61 = ptr + 1'h1; // @[WriteMemoryController.scala 146:18]
  assign _GEN_14 = _T_58 ? {{7'd0}, _T_59} : _GEN_10; // @[WriteMemoryController.scala 142:29]
  assign _GEN_18 = _T_57 ? _GEN_14 : _GEN_10; // @[WriteMemoryController.scala 139:76]
  assign _T_62 = state == 2'h2; // @[WriteMemoryController.scala 156:15]
  assign _T_64 = _T_62 & io_MemResp_valid; // @[WriteMemoryController.scala 156:32]
  assign _T_65 = sendbytemask == 8'h0; // @[WriteMemoryController.scala 158:27]
  assign _T_68 = io_output_ready & io_output_valid; // @[Decoupled.scala 40:37]
  assign io_NodeReq_ready = state == 2'h0; // @[WriteMemoryController.scala 87:20]
  assign io_MemReq_valid = _T_55 & _T_56; // @[WriteMemoryController.scala 99:19 WriteMemoryController.scala 140:21]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_29; // @[WriteMemoryController.scala 100:23]
  assign io_MemReq_bits_data = ptr ? linebuffer_1 : linebuffer_0; // @[WriteMemoryController.scala 102:23]
  assign io_MemReq_bits_mask = sendbytemask[3:0]; // @[WriteMemoryController.scala 103:23]
  assign io_MemReq_bits_tag = {{7'd0}, myID}; // @[WriteMemoryController.scala 107:22]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[WriteMemoryController.scala 110:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[WriteMemoryController.scala 109:26]
  assign io_output_valid = state == 2'h3; // @[WriteMemoryController.scala 95:19 WriteMemoryController.scala 168:21]
  assign io_free = state == 2'h0; // @[WriteMemoryController.scala 85:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ID = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sendbytemask = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ReqAddress = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ptr = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  linebuffer_0 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  linebuffer_1 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  myID = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  isWrite = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    ID <= reset | ID;
    if (reset) begin
      request_R_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_18[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_9) begin
        ReqAddress <= {{10'd0}, _T_11};
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (_T_4) begin
        ptr <= 1'h0;
      end else begin
        if (_T_57) begin
          if (_T_58) begin
            ptr <= _T_61;
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (_T_9) begin
        linebuffer_0 <= _T_53;
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (_T_9) begin
        linebuffer_1 <= _T_54;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_4) begin
        if (_T_68) begin
          state <= 2'h0;
        end else begin
          if (_T_64) begin
            if (_T_65) begin
              state <= 2'h3;
            end else begin
              state <= 2'h1;
            end
          end else begin
            if (_T_57) begin
              if (_T_58) begin
                state <= 2'h2;
              end else begin
                if (_T_9) begin
                  state <= 2'h1;
                end
              end
            end else begin
              if (_T_9) begin
                state <= 2'h1;
              end
            end
          end
        end
      end else begin
        if (_T_64) begin
          if (_T_65) begin
            state <= 2'h3;
          end else begin
            state <= 2'h1;
          end
        end else begin
          if (_T_57) begin
            if (_T_58) begin
              state <= 2'h2;
            end else begin
              if (_T_9) begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_9) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      myID <= 1'h0;
    end else begin
      myID <= ID;
    end
    if (reset) begin
      isWrite <= 1'h0;
    end else begin
      isWrite <= 1'h1;
    end
  end
endmodule
module WriteMemoryController(
  input         clock,
  input         reset,
  output        io_WriteIn_0_ready,
  input         io_WriteIn_0_valid,
  input  [21:0] io_WriteIn_0_bits_address,
  input  [31:0] io_WriteIn_0_bits_data,
  input  [4:0]  io_WriteIn_0_bits_taskID,
  output        io_WriteOut_0_valid,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag
);
  wire  in_arb_io_in_0_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_0_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_0_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_0_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_0_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_out_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_out_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_out_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_out_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire [7:0] in_arb_io_out_bits_Typ; // @[WriteMemoryController.scala 194:25]
  wire  alloc_arb_io_in_0_ready; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_in_0_valid; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_in_1_ready; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_in_1_valid; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_out_ready; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_out_valid; // @[WriteMemoryController.scala 196:25]
  wire  cachereq_arb_io_in_0_ready; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_0_valid; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_0_bits_addr; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_0_bits_data; // @[WriteMemoryController.scala 199:31]
  wire [3:0] cachereq_arb_io_in_0_bits_mask; // @[WriteMemoryController.scala 199:31]
  wire [7:0] cachereq_arb_io_in_0_bits_tag; // @[WriteMemoryController.scala 199:31]
  wire [4:0] cachereq_arb_io_in_0_bits_taskID; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_0_bits_iswrite; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_1_ready; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_1_valid; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_1_bits_addr; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_1_bits_data; // @[WriteMemoryController.scala 199:31]
  wire [3:0] cachereq_arb_io_in_1_bits_mask; // @[WriteMemoryController.scala 199:31]
  wire [7:0] cachereq_arb_io_in_1_bits_tag; // @[WriteMemoryController.scala 199:31]
  wire [4:0] cachereq_arb_io_in_1_bits_taskID; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_1_bits_iswrite; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_out_ready; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_out_valid; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_out_bits_addr; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_out_bits_data; // @[WriteMemoryController.scala 199:31]
  wire [3:0] cachereq_arb_io_out_bits_mask; // @[WriteMemoryController.scala 199:31]
  wire [7:0] cachereq_arb_io_out_bits_tag; // @[WriteMemoryController.scala 199:31]
  wire [4:0] cachereq_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_out_bits_iswrite; // @[WriteMemoryController.scala 199:31]
  wire  cacheresp_demux_io_en; // @[WriteMemoryController.scala 201:31]
  wire [31:0] cacheresp_demux_io_input_data; // @[WriteMemoryController.scala 201:31]
  wire [7:0] cacheresp_demux_io_input_tag; // @[WriteMemoryController.scala 201:31]
  wire  cacheresp_demux_io_sel; // @[WriteMemoryController.scala 201:31]
  wire  cacheresp_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 201:31]
  wire [31:0] cacheresp_demux_io_outputs_0_data; // @[WriteMemoryController.scala 201:31]
  wire [7:0] cacheresp_demux_io_outputs_0_tag; // @[WriteMemoryController.scala 201:31]
  wire  cacheresp_demux_io_outputs_1_valid; // @[WriteMemoryController.scala 201:31]
  wire [31:0] cacheresp_demux_io_outputs_1_data; // @[WriteMemoryController.scala 201:31]
  wire [7:0] cacheresp_demux_io_outputs_1_tag; // @[WriteMemoryController.scala 201:31]
  wire  out_arb_clock; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_0_ready; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_0_valid; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_1_ready; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_1_valid; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_out_ready; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_out_valid; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_chosen; // @[WriteMemoryController.scala 204:25]
  wire  out_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_enable; // @[WriteMemoryController.scala 205:25]
  wire  WriteTable_0_clock; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_reset; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_NodeReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_NodeReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [21:0] WriteTable_0_io_NodeReq_bits_address; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_0_io_NodeReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [4:0] WriteTable_0_io_NodeReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire [7:0] WriteTable_0_io_NodeReq_bits_Typ; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_0_io_MemReq_bits_addr; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_0_io_MemReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [3:0] WriteTable_0_io_MemReq_bits_mask; // @[WriteMemoryController.scala 223:29]
  wire [4:0] WriteTable_0_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemResp_valid; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_output_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_output_valid; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_free; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_clock; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_reset; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_NodeReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_NodeReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [21:0] WriteTable_1_io_NodeReq_bits_address; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_1_io_NodeReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [4:0] WriteTable_1_io_NodeReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire [7:0] WriteTable_1_io_NodeReq_bits_Typ; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_1_io_MemReq_bits_addr; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_1_io_MemReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [3:0] WriteTable_1_io_MemReq_bits_mask; // @[WriteMemoryController.scala 223:29]
  wire [7:0] WriteTable_1_io_MemReq_bits_tag; // @[WriteMemoryController.scala 223:29]
  wire [4:0] WriteTable_1_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemResp_valid; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_output_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_output_valid; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_free; // @[WriteMemoryController.scala 223:29]
  ArbiterTree in_arb ( // @[WriteMemoryController.scala 194:25]
    .io_in_0_ready(in_arb_io_in_0_ready),
    .io_in_0_valid(in_arb_io_in_0_valid),
    .io_in_0_bits_address(in_arb_io_in_0_bits_address),
    .io_in_0_bits_data(in_arb_io_in_0_bits_data),
    .io_in_0_bits_taskID(in_arb_io_in_0_bits_taskID),
    .io_out_ready(in_arb_io_out_ready),
    .io_out_valid(in_arb_io_out_valid),
    .io_out_bits_address(in_arb_io_out_bits_address),
    .io_out_bits_data(in_arb_io_out_bits_data),
    .io_out_bits_taskID(in_arb_io_out_bits_taskID),
    .io_out_bits_Typ(in_arb_io_out_bits_Typ)
  );
  Arbiter alloc_arb ( // @[WriteMemoryController.scala 196:25]
    .io_in_0_ready(alloc_arb_io_in_0_ready),
    .io_in_0_valid(alloc_arb_io_in_0_valid),
    .io_in_1_ready(alloc_arb_io_in_1_ready),
    .io_in_1_valid(alloc_arb_io_in_1_valid),
    .io_out_ready(alloc_arb_io_out_ready),
    .io_out_valid(alloc_arb_io_out_valid)
  );
  Arbiter_1 cachereq_arb ( // @[WriteMemoryController.scala 199:31]
    .io_in_0_ready(cachereq_arb_io_in_0_ready),
    .io_in_0_valid(cachereq_arb_io_in_0_valid),
    .io_in_0_bits_addr(cachereq_arb_io_in_0_bits_addr),
    .io_in_0_bits_data(cachereq_arb_io_in_0_bits_data),
    .io_in_0_bits_mask(cachereq_arb_io_in_0_bits_mask),
    .io_in_0_bits_tag(cachereq_arb_io_in_0_bits_tag),
    .io_in_0_bits_taskID(cachereq_arb_io_in_0_bits_taskID),
    .io_in_0_bits_iswrite(cachereq_arb_io_in_0_bits_iswrite),
    .io_in_1_ready(cachereq_arb_io_in_1_ready),
    .io_in_1_valid(cachereq_arb_io_in_1_valid),
    .io_in_1_bits_addr(cachereq_arb_io_in_1_bits_addr),
    .io_in_1_bits_data(cachereq_arb_io_in_1_bits_data),
    .io_in_1_bits_mask(cachereq_arb_io_in_1_bits_mask),
    .io_in_1_bits_tag(cachereq_arb_io_in_1_bits_tag),
    .io_in_1_bits_taskID(cachereq_arb_io_in_1_bits_taskID),
    .io_in_1_bits_iswrite(cachereq_arb_io_in_1_bits_iswrite),
    .io_out_ready(cachereq_arb_io_out_ready),
    .io_out_valid(cachereq_arb_io_out_valid),
    .io_out_bits_addr(cachereq_arb_io_out_bits_addr),
    .io_out_bits_data(cachereq_arb_io_out_bits_data),
    .io_out_bits_mask(cachereq_arb_io_out_bits_mask),
    .io_out_bits_tag(cachereq_arb_io_out_bits_tag),
    .io_out_bits_taskID(cachereq_arb_io_out_bits_taskID),
    .io_out_bits_iswrite(cachereq_arb_io_out_bits_iswrite)
  );
  Demux cacheresp_demux ( // @[WriteMemoryController.scala 201:31]
    .io_en(cacheresp_demux_io_en),
    .io_input_data(cacheresp_demux_io_input_data),
    .io_input_tag(cacheresp_demux_io_input_tag),
    .io_sel(cacheresp_demux_io_sel),
    .io_outputs_0_valid(cacheresp_demux_io_outputs_0_valid),
    .io_outputs_0_data(cacheresp_demux_io_outputs_0_data),
    .io_outputs_0_tag(cacheresp_demux_io_outputs_0_tag),
    .io_outputs_1_valid(cacheresp_demux_io_outputs_1_valid),
    .io_outputs_1_data(cacheresp_demux_io_outputs_1_data),
    .io_outputs_1_tag(cacheresp_demux_io_outputs_1_tag)
  );
  RRArbiter out_arb ( // @[WriteMemoryController.scala 204:25]
    .clock(out_arb_clock),
    .io_in_0_ready(out_arb_io_in_0_ready),
    .io_in_0_valid(out_arb_io_in_0_valid),
    .io_in_1_ready(out_arb_io_in_1_ready),
    .io_in_1_valid(out_arb_io_in_1_valid),
    .io_out_ready(out_arb_io_out_ready),
    .io_out_valid(out_arb_io_out_valid),
    .io_chosen(out_arb_io_chosen)
  );
  DeMuxTree out_demux ( // @[WriteMemoryController.scala 205:25]
    .io_outputs_0_valid(out_demux_io_outputs_0_valid),
    .io_enable(out_demux_io_enable)
  );
  WriteTableEntry WriteTable_0 ( // @[WriteMemoryController.scala 223:29]
    .clock(WriteTable_0_clock),
    .reset(WriteTable_0_reset),
    .io_NodeReq_ready(WriteTable_0_io_NodeReq_ready),
    .io_NodeReq_valid(WriteTable_0_io_NodeReq_valid),
    .io_NodeReq_bits_address(WriteTable_0_io_NodeReq_bits_address),
    .io_NodeReq_bits_data(WriteTable_0_io_NodeReq_bits_data),
    .io_NodeReq_bits_taskID(WriteTable_0_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(WriteTable_0_io_NodeReq_bits_Typ),
    .io_MemReq_ready(WriteTable_0_io_MemReq_ready),
    .io_MemReq_valid(WriteTable_0_io_MemReq_valid),
    .io_MemReq_bits_addr(WriteTable_0_io_MemReq_bits_addr),
    .io_MemReq_bits_data(WriteTable_0_io_MemReq_bits_data),
    .io_MemReq_bits_mask(WriteTable_0_io_MemReq_bits_mask),
    .io_MemReq_bits_taskID(WriteTable_0_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(WriteTable_0_io_MemReq_bits_iswrite),
    .io_MemResp_valid(WriteTable_0_io_MemResp_valid),
    .io_output_ready(WriteTable_0_io_output_ready),
    .io_output_valid(WriteTable_0_io_output_valid),
    .io_free(WriteTable_0_io_free)
  );
  WriteTableEntry_1 WriteTable_1 ( // @[WriteMemoryController.scala 223:29]
    .clock(WriteTable_1_clock),
    .reset(WriteTable_1_reset),
    .io_NodeReq_ready(WriteTable_1_io_NodeReq_ready),
    .io_NodeReq_valid(WriteTable_1_io_NodeReq_valid),
    .io_NodeReq_bits_address(WriteTable_1_io_NodeReq_bits_address),
    .io_NodeReq_bits_data(WriteTable_1_io_NodeReq_bits_data),
    .io_NodeReq_bits_taskID(WriteTable_1_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(WriteTable_1_io_NodeReq_bits_Typ),
    .io_MemReq_ready(WriteTable_1_io_MemReq_ready),
    .io_MemReq_valid(WriteTable_1_io_MemReq_valid),
    .io_MemReq_bits_addr(WriteTable_1_io_MemReq_bits_addr),
    .io_MemReq_bits_data(WriteTable_1_io_MemReq_bits_data),
    .io_MemReq_bits_mask(WriteTable_1_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(WriteTable_1_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(WriteTable_1_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(WriteTable_1_io_MemReq_bits_iswrite),
    .io_MemResp_valid(WriteTable_1_io_MemResp_valid),
    .io_output_ready(WriteTable_1_io_output_ready),
    .io_output_valid(WriteTable_1_io_output_valid),
    .io_free(WriteTable_1_io_free)
  );
  assign io_WriteIn_0_ready = in_arb_io_in_0_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteOut_0_valid = out_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 214:20]
  assign io_MemReq_valid = cachereq_arb_io_out_valid; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_addr = cachereq_arb_io_out_bits_addr; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_data = cachereq_arb_io_out_bits_data; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_mask = cachereq_arb_io_out_bits_mask; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_tag = cachereq_arb_io_out_bits_tag; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_taskID = cachereq_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_iswrite = cachereq_arb_io_out_bits_iswrite; // @[WriteMemoryController.scala 261:13]
  assign in_arb_io_in_0_valid = io_WriteIn_0_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_0_bits_address = io_WriteIn_0_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_0_bits_data = io_WriteIn_0_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_0_bits_taskID = io_WriteIn_0_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_out_ready = alloc_arb_io_out_valid; // @[WriteMemoryController.scala 256:23]
  assign alloc_arb_io_in_0_valid = WriteTable_0_io_free; // @[WriteMemoryController.scala 226:30]
  assign alloc_arb_io_in_1_valid = WriteTable_1_io_free; // @[WriteMemoryController.scala 226:30]
  assign alloc_arb_io_out_ready = in_arb_io_out_valid; // @[WriteMemoryController.scala 257:26]
  assign cachereq_arb_io_in_0_valid = WriteTable_0_io_MemReq_valid; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_addr = WriteTable_0_io_MemReq_bits_addr; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_data = WriteTable_0_io_MemReq_bits_data; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_mask = WriteTable_0_io_MemReq_bits_mask; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_tag = 8'h0; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_taskID = WriteTable_0_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_iswrite = WriteTable_0_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_valid = WriteTable_1_io_MemReq_valid; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_addr = WriteTable_1_io_MemReq_bits_addr; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_data = WriteTable_1_io_MemReq_bits_data; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_mask = WriteTable_1_io_MemReq_bits_mask; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_tag = WriteTable_1_io_MemReq_bits_tag; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_taskID = WriteTable_1_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_iswrite = WriteTable_1_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_out_ready = io_MemReq_ready; // @[WriteMemoryController.scala 261:13]
  assign cacheresp_demux_io_en = io_MemResp_valid; // @[WriteMemoryController.scala 264:25]
  assign cacheresp_demux_io_input_data = io_MemResp_bits_data; // @[WriteMemoryController.scala 265:28]
  assign cacheresp_demux_io_input_tag = io_MemResp_bits_tag; // @[WriteMemoryController.scala 265:28]
  assign cacheresp_demux_io_sel = io_MemResp_bits_tag[0]; // @[WriteMemoryController.scala 266:26]
  assign out_arb_clock = clock;
  assign out_arb_io_in_0_valid = WriteTable_0_io_output_valid; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_in_1_valid = WriteTable_1_io_output_valid; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_out_ready = 1'h1; // @[WriteMemoryController.scala 269:24]
  assign out_demux_io_enable = out_arb_io_out_ready & out_arb_io_out_valid; // @[WriteMemoryController.scala 270:23]
  assign WriteTable_0_clock = clock;
  assign WriteTable_0_reset = reset;
  assign WriteTable_0_io_NodeReq_valid = alloc_arb_io_in_0_ready & alloc_arb_io_in_0_valid; // @[WriteMemoryController.scala 228:34]
  assign WriteTable_0_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_data = in_arb_io_out_bits_data; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_MemReq_ready = cachereq_arb_io_in_0_ready; // @[WriteMemoryController.scala 232:27]
  assign WriteTable_0_io_MemResp_valid = cacheresp_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 235:28]
  assign WriteTable_0_io_output_ready = out_arb_io_in_0_ready; // @[WriteMemoryController.scala 238:22]
  assign WriteTable_1_clock = clock;
  assign WriteTable_1_reset = reset;
  assign WriteTable_1_io_NodeReq_valid = alloc_arb_io_in_1_ready & alloc_arb_io_in_1_valid; // @[WriteMemoryController.scala 228:34]
  assign WriteTable_1_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_data = in_arb_io_out_bits_data; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_MemReq_ready = cachereq_arb_io_in_1_ready; // @[WriteMemoryController.scala 232:27]
  assign WriteTable_1_io_MemResp_valid = cacheresp_demux_io_outputs_1_valid; // @[WriteMemoryController.scala 235:28]
  assign WriteTable_1_io_output_ready = out_arb_io_in_1_ready; // @[WriteMemoryController.scala 238:22]
endmodule
module LockingRRArbiter_1(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_address,
  input  [4:0]  io_in_0_bits_taskID,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_address,
  input  [4:0]  io_in_1_bits_taskID,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [31:0] io_out_bits_address,
  output [4:0]  io_out_bits_taskID,
  output        io_chosen
);
  wire  _T; // @[Decoupled.scala 40:37]
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Arbiter.scala 67:57]
  wire  _T_5; // @[Arbiter.scala 68:83]
  wire  _T_7; // @[Arbiter.scala 31:68]
  wire  _T_9; // @[Arbiter.scala 31:78]
  wire  _T_10; // @[Arbiter.scala 31:78]
  wire  _T_14; // @[Arbiter.scala 72:50]
  wire  _GEN_13; // @[Arbiter.scala 77:27]
  assign _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = 1'h1 > _T_1; // @[Arbiter.scala 67:57]
  assign _T_5 = io_in_1_valid & _T_3; // @[Arbiter.scala 68:83]
  assign _T_7 = _T_5 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_9 = _T_5 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_10 = _T_7 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_14 = _T_3 | _T_10; // @[Arbiter.scala 72:50]
  assign _GEN_13 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_9 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_14 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_RouteID = io_chosen ? 16'h1 : 16'h0; // @[Arbiter.scala 42:15]
  assign io_out_bits_address = io_chosen ? io_in_1_bits_address : io_in_0_bits_address; // @[Arbiter.scala 42:15]
  assign io_out_bits_taskID = io_chosen ? io_in_1_bits_taskID : io_in_0_bits_taskID; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_5 | _GEN_13; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (_T) begin
      _T_1 <= io_chosen;
    end
  end
endmodule
module ArbiterTree_1(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_address,
  input  [4:0]  io_in_0_bits_taskID,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_address,
  input  [4:0]  io_in_1_bits_taskID,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [31:0] io_out_bits_address,
  output [4:0]  io_out_bits_taskID
);
  wire  LockingRRArbiter_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_chosen; // @[ArbiterTree.scala 32:13]
  LockingRRArbiter_1 LockingRRArbiter ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_clock),
    .io_in_0_ready(LockingRRArbiter_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_io_in_0_valid),
    .io_in_0_bits_address(LockingRRArbiter_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_io_in_0_bits_taskID),
    .io_in_1_ready(LockingRRArbiter_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_io_in_1_valid),
    .io_in_1_bits_address(LockingRRArbiter_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_io_in_1_bits_taskID),
    .io_out_ready(LockingRRArbiter_io_out_ready),
    .io_out_valid(LockingRRArbiter_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_io_out_bits_taskID),
    .io_chosen(LockingRRArbiter_io_chosen)
  );
  assign io_in_0_ready = LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_1_ready = LockingRRArbiter_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_out_valid = LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_RouteID = LockingRRArbiter_io_out_bits_RouteID; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_address = LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_taskID = LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 65:12]
  assign LockingRRArbiter_clock = clock;
  assign LockingRRArbiter_io_in_0_valid = io_in_0_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_address = io_in_0_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_taskID = io_in_0_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_valid = io_in_1_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_address = io_in_1_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_taskID = io_in_1_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_out_ready = io_out_ready; // @[ArbiterTree.scala 65:12]
endmodule
module RRArbiter_1(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [15:0] io_in_0_bits_RouteID,
  input  [31:0] io_in_0_bits_data,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [15:0] io_in_1_bits_RouteID,
  input  [31:0] io_in_1_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [31:0] io_out_bits_data,
  output        io_chosen
);
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Arbiter.scala 67:57]
  wire  _T_5; // @[Arbiter.scala 68:83]
  wire  _T_7; // @[Arbiter.scala 31:68]
  wire  _T_10; // @[Arbiter.scala 31:78]
  wire  _GEN_11; // @[Arbiter.scala 77:27]
  assign _T_3 = 1'h1 > _T_1; // @[Arbiter.scala 67:57]
  assign _T_5 = io_in_1_valid & _T_3; // @[Arbiter.scala 68:83]
  assign _T_7 = _T_5 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_10 = _T_7 == 1'h0; // @[Arbiter.scala 31:78]
  assign _GEN_11 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_5 == 1'h0; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_3 | _T_10; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_RouteID = io_chosen ? io_in_1_bits_RouteID : io_in_0_bits_RouteID; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_5 | _GEN_11; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_out_valid) begin
      _T_1 <= io_chosen;
    end
  end
endmodule
module Demux_3(
  input         io_en,
  input  [31:0] io_input_data,
  input         io_sel,
  output        io_outputs_0_valid,
  output [31:0] io_outputs_0_data,
  output        io_outputs_1_valid,
  output [31:0] io_outputs_1_data
);
  wire  _GEN_0; // @[Muxes.scala 29:25]
  assign _GEN_0 = 1'h0 == io_sel; // @[Muxes.scala 29:25]
  assign io_outputs_0_valid = io_en & _GEN_0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_0_data = io_input_data; // @[Muxes.scala 23:19]
  assign io_outputs_1_valid = io_en & io_sel; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_1_data = io_input_data; // @[Muxes.scala 23:19]
endmodule
module DeMuxTree_1(
  output        io_outputs_0_valid,
  output [31:0] io_outputs_0_data,
  output        io_outputs_1_valid,
  output [31:0] io_outputs_1_data,
  input  [15:0] io_input_RouteID,
  input  [31:0] io_input_data,
  input         io_enable
);
  wire  Demux_io_en; // @[Muxes.scala 91:13]
  wire [31:0] Demux_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [31:0] Demux_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [31:0] Demux_io_outputs_1_data; // @[Muxes.scala 91:13]
  Demux_3 Demux ( // @[Muxes.scala 91:13]
    .io_en(Demux_io_en),
    .io_input_data(Demux_io_input_data),
    .io_sel(Demux_io_sel),
    .io_outputs_0_valid(Demux_io_outputs_0_valid),
    .io_outputs_0_data(Demux_io_outputs_0_data),
    .io_outputs_1_valid(Demux_io_outputs_1_valid),
    .io_outputs_1_data(Demux_io_outputs_1_data)
  );
  assign io_outputs_0_valid = Demux_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_0_data = Demux_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_1_valid = Demux_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_1_data = Demux_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign Demux_io_en = io_enable; // @[Muxes.scala 135:14]
  assign Demux_io_input_data = io_input_data; // @[Muxes.scala 134:17]
  assign Demux_io_sel = io_input_RouteID[0]; // @[Muxes.scala 136:15]
endmodule
module ReadTableEntry(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [15:0] io_NodeReq_bits_RouteID,
  input  [31:0] io_NodeReq_bits_address,
  input  [4:0]  io_NodeReq_bits_taskID,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_data,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output [31:0] io_output_bits_data,
  output        io_free
);
  reg  ID; // @[ReadMemoryController.scala 49:19]
  reg [31:0] _RAND_0;
  reg [15:0] request_R_RouteID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_1;
  reg [31:0] request_R_address; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_2;
  reg [4:0] request_R_taskID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_3;
  reg [63:0] bitmask; // @[ReadMemoryController.scala 56:29]
  reg [63:0] _RAND_4;
  reg [7:0] sendbytemask; // @[ReadMemoryController.scala 58:29]
  reg [31:0] _RAND_5;
  reg [31:0] ReqAddress; // @[ReadMemoryController.scala 62:27]
  reg [31:0] _RAND_6;
  reg  ptr; // @[ReadMemoryController.scala 66:27]
  reg [31:0] _RAND_7;
  reg [31:0] linebuffer_0; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_8;
  reg [31:0] linebuffer_1; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[ReadMemoryController.scala 73:68]
  reg [31:0] _RAND_10;
  wire [2:0] _T_6; // @[Cat.scala 29:58]
  wire [31:0] _GEN_57; // @[ReadMemoryController.scala 96:37]
  reg  isWrite; // @[ReadMemoryController.scala 100:24]
  reg [31:0] _RAND_11;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire [29:0] _T_10; // @[ReadMemoryController.scala 115:44]
  wire [31:0] _T_11; // @[ReadMemoryController.scala 115:69]
  wire [1:0] _T_28; // @[helpers.scala 39:32]
  wire [4:0] _T_29; // @[Cat.scala 29:58]
  wire [94:0] _T_30; // @[helpers.scala 40:26]
  wire [10:0] _T_47; // @[helpers.scala 20:26]
  wire [94:0] _GEN_5; // @[ReadMemoryController.scala 111:28]
  wire [10:0] _GEN_6; // @[ReadMemoryController.scala 111:28]
  wire  _T_48; // @[Conditional.scala 37:30]
  wire  _T_50; // @[Conditional.scala 37:30]
  wire [3:0] _T_51; // @[ReadMemoryController.scala 144:38]
  wire [10:0] _GEN_8; // @[ReadMemoryController.scala 142:29]
  wire  _T_52; // @[Conditional.scala 37:30]
  wire  _T_54; // @[ReadMemoryController.scala 154:20]
  wire  _T_55; // @[ReadMemoryController.scala 156:27]
  wire  _T_56; // @[Conditional.scala 37:30]
  wire [63:0] _T_57; // @[ReadMemoryController.scala 165:29]
  wire [63:0] _T_58; // @[ReadMemoryController.scala 165:36]
  wire [1:0] _T_59; // @[ReadMemoryController.scala 165:71]
  wire [4:0] _T_60; // @[Cat.scala 29:58]
  wire [63:0] _T_61; // @[ReadMemoryController.scala 165:47]
  wire [63:0] _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_31; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_42; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_53; // @[Conditional.scala 40:58]
  wire [31:0] output_; // @[ReadMemoryController.scala 165:14]
  wire [31:0] _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_43; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_48; // @[Conditional.scala 40:58]
  assign _T_6 = {ptr,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_57 = {{29'd0}, _T_6}; // @[ReadMemoryController.scala 96:37]
  assign _T_9 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_NodeReq_bits_address[31:2]; // @[ReadMemoryController.scala 115:44]
  assign _T_11 = {_T_10, 2'h0}; // @[ReadMemoryController.scala 115:69]
  assign _T_28 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_29 = {_T_28,3'h0}; // @[Cat.scala 29:58]
  assign _T_30 = 95'hffffffff << _T_29; // @[helpers.scala 40:26]
  assign _T_47 = 11'hf << _T_28; // @[helpers.scala 20:26]
  assign _GEN_5 = _T_9 ? _T_30 : {{31'd0}, bitmask}; // @[ReadMemoryController.scala 111:28]
  assign _GEN_6 = _T_9 ? _T_47 : {{3'd0}, sendbytemask}; // @[ReadMemoryController.scala 111:28]
  assign _T_48 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_50 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_51 = sendbytemask[7:4]; // @[ReadMemoryController.scala 144:38]
  assign _GEN_8 = io_MemReq_ready ? {{7'd0}, _T_51} : _GEN_6; // @[ReadMemoryController.scala 142:29]
  assign _T_52 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_54 = ptr + 1'h1; // @[ReadMemoryController.scala 154:20]
  assign _T_55 = sendbytemask == 8'h0; // @[ReadMemoryController.scala 156:27]
  assign _T_56 = 2'h3 == state; // @[Conditional.scala 37:30]
  assign _T_57 = {linebuffer_1,linebuffer_0}; // @[ReadMemoryController.scala 165:29]
  assign _T_58 = _T_57 & bitmask; // @[ReadMemoryController.scala 165:36]
  assign _T_59 = request_R_address[1:0]; // @[ReadMemoryController.scala 165:71]
  assign _T_60 = {_T_59,3'h0}; // @[Cat.scala 29:58]
  assign _T_61 = _T_58 >> _T_60; // @[ReadMemoryController.scala 165:47]
  assign _GEN_20 = _T_56 ? _T_61 : 64'h0; // @[Conditional.scala 39:67]
  assign _GEN_31 = _T_52 ? 64'h0 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_50 ? 64'h0 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_53 = _T_48 ? 64'h0 : _GEN_42; // @[Conditional.scala 40:58]
  assign output_ = _GEN_53[31:0]; // @[ReadMemoryController.scala 165:14]
  assign _GEN_21 = _T_56 ? output_ : 32'h0; // @[Conditional.scala 39:67]
  assign _GEN_30 = _T_52 ? 1'h0 : _T_56; // @[Conditional.scala 39:67]
  assign _GEN_32 = _T_52 ? 32'h0 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_50 ? _GEN_8 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_41 = _T_50 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_43 = _T_50 ? 32'h0 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_48 = _T_48 ? _GEN_6 : _GEN_36; // @[Conditional.scala 40:58]
  assign io_NodeReq_ready = state == 2'h0; // @[ReadMemoryController.scala 83:20]
  assign io_MemReq_valid = _T_48 ? 1'h0 : _T_50; // @[ReadMemoryController.scala 95:19 ReadMemoryController.scala 140:23]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_57; // @[ReadMemoryController.scala 96:23]
  assign io_MemReq_bits_tag = {{7'd0}, ID}; // @[ReadMemoryController.scala 99:22]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[ReadMemoryController.scala 104:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[ReadMemoryController.scala 101:26]
  assign io_output_valid = _T_48 ? 1'h0 : _GEN_41; // @[ReadMemoryController.scala 90:19 ReadMemoryController.scala 164:23]
  assign io_output_bits_RouteID = request_R_RouteID; // @[ReadMemoryController.scala 91:26]
  assign io_output_bits_data = _T_48 ? 32'h0 : _GEN_43; // @[ReadMemoryController.scala 93:23 ReadMemoryController.scala 168:29]
  assign io_free = state == 2'h0; // @[ReadMemoryController.scala 81:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ID = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_RouteID = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  request_R_address = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  request_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  bitmask = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sendbytemask = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ReqAddress = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ptr = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  linebuffer_0 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  linebuffer_1 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  isWrite = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    ID <= reset;
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_9) begin
        request_R_RouteID <= io_NodeReq_bits_RouteID;
      end
    end
    if (reset) begin
      request_R_address <= 32'h0;
    end else begin
      if (_T_9) begin
        request_R_address <= io_NodeReq_bits_address;
      end
    end
    if (reset) begin
      request_R_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      bitmask <= 64'h0;
    end else begin
      bitmask <= _GEN_5[63:0];
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_48[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_9) begin
        ReqAddress <= _T_11;
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              ptr <= _T_54;
            end
          end else begin
            if (_T_56) begin
              ptr <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (1'h0 == ptr) begin
                linebuffer_0 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (ptr) begin
                linebuffer_1 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_48) begin
        if (_T_9) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_50) begin
          if (io_MemReq_ready) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (_T_55) begin
                state <= 2'h3;
              end else begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_56) begin
              if (io_output_ready) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    isWrite <= reset;
  end
endmodule
module ReadTableEntry_1(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [15:0] io_NodeReq_bits_RouteID,
  input  [31:0] io_NodeReq_bits_address,
  input  [4:0]  io_NodeReq_bits_taskID,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_data,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output [31:0] io_output_bits_data,
  output        io_free
);
  reg  ID; // @[ReadMemoryController.scala 49:19]
  reg [31:0] _RAND_0;
  reg [15:0] request_R_RouteID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_1;
  reg [31:0] request_R_address; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_2;
  reg [4:0] request_R_taskID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_3;
  reg [63:0] bitmask; // @[ReadMemoryController.scala 56:29]
  reg [63:0] _RAND_4;
  reg [7:0] sendbytemask; // @[ReadMemoryController.scala 58:29]
  reg [31:0] _RAND_5;
  reg [31:0] ReqAddress; // @[ReadMemoryController.scala 62:27]
  reg [31:0] _RAND_6;
  reg  ptr; // @[ReadMemoryController.scala 66:27]
  reg [31:0] _RAND_7;
  reg [31:0] linebuffer_0; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_8;
  reg [31:0] linebuffer_1; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[ReadMemoryController.scala 73:68]
  reg [31:0] _RAND_10;
  wire [2:0] _T_6; // @[Cat.scala 29:58]
  wire [31:0] _GEN_57; // @[ReadMemoryController.scala 96:37]
  reg  isWrite; // @[ReadMemoryController.scala 100:24]
  reg [31:0] _RAND_11;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire [29:0] _T_10; // @[ReadMemoryController.scala 115:44]
  wire [31:0] _T_11; // @[ReadMemoryController.scala 115:69]
  wire [1:0] _T_28; // @[helpers.scala 39:32]
  wire [4:0] _T_29; // @[Cat.scala 29:58]
  wire [94:0] _T_30; // @[helpers.scala 40:26]
  wire [10:0] _T_47; // @[helpers.scala 20:26]
  wire [94:0] _GEN_5; // @[ReadMemoryController.scala 111:28]
  wire [10:0] _GEN_6; // @[ReadMemoryController.scala 111:28]
  wire  _T_48; // @[Conditional.scala 37:30]
  wire  _T_50; // @[Conditional.scala 37:30]
  wire [3:0] _T_51; // @[ReadMemoryController.scala 144:38]
  wire [10:0] _GEN_8; // @[ReadMemoryController.scala 142:29]
  wire  _T_52; // @[Conditional.scala 37:30]
  wire  _T_54; // @[ReadMemoryController.scala 154:20]
  wire  _T_55; // @[ReadMemoryController.scala 156:27]
  wire  _T_56; // @[Conditional.scala 37:30]
  wire [63:0] _T_57; // @[ReadMemoryController.scala 165:29]
  wire [63:0] _T_58; // @[ReadMemoryController.scala 165:36]
  wire [1:0] _T_59; // @[ReadMemoryController.scala 165:71]
  wire [4:0] _T_60; // @[Cat.scala 29:58]
  wire [63:0] _T_61; // @[ReadMemoryController.scala 165:47]
  wire [63:0] _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_31; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_42; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_53; // @[Conditional.scala 40:58]
  wire [31:0] output_; // @[ReadMemoryController.scala 165:14]
  wire [31:0] _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_43; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_48; // @[Conditional.scala 40:58]
  assign _T_6 = {ptr,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_57 = {{29'd0}, _T_6}; // @[ReadMemoryController.scala 96:37]
  assign _T_9 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_NodeReq_bits_address[31:2]; // @[ReadMemoryController.scala 115:44]
  assign _T_11 = {_T_10, 2'h0}; // @[ReadMemoryController.scala 115:69]
  assign _T_28 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_29 = {_T_28,3'h0}; // @[Cat.scala 29:58]
  assign _T_30 = 95'hffffffff << _T_29; // @[helpers.scala 40:26]
  assign _T_47 = 11'hf << _T_28; // @[helpers.scala 20:26]
  assign _GEN_5 = _T_9 ? _T_30 : {{31'd0}, bitmask}; // @[ReadMemoryController.scala 111:28]
  assign _GEN_6 = _T_9 ? _T_47 : {{3'd0}, sendbytemask}; // @[ReadMemoryController.scala 111:28]
  assign _T_48 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_50 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_51 = sendbytemask[7:4]; // @[ReadMemoryController.scala 144:38]
  assign _GEN_8 = io_MemReq_ready ? {{7'd0}, _T_51} : _GEN_6; // @[ReadMemoryController.scala 142:29]
  assign _T_52 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_54 = ptr + 1'h1; // @[ReadMemoryController.scala 154:20]
  assign _T_55 = sendbytemask == 8'h0; // @[ReadMemoryController.scala 156:27]
  assign _T_56 = 2'h3 == state; // @[Conditional.scala 37:30]
  assign _T_57 = {linebuffer_1,linebuffer_0}; // @[ReadMemoryController.scala 165:29]
  assign _T_58 = _T_57 & bitmask; // @[ReadMemoryController.scala 165:36]
  assign _T_59 = request_R_address[1:0]; // @[ReadMemoryController.scala 165:71]
  assign _T_60 = {_T_59,3'h0}; // @[Cat.scala 29:58]
  assign _T_61 = _T_58 >> _T_60; // @[ReadMemoryController.scala 165:47]
  assign _GEN_20 = _T_56 ? _T_61 : 64'h0; // @[Conditional.scala 39:67]
  assign _GEN_31 = _T_52 ? 64'h0 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_50 ? 64'h0 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_53 = _T_48 ? 64'h0 : _GEN_42; // @[Conditional.scala 40:58]
  assign output_ = _GEN_53[31:0]; // @[ReadMemoryController.scala 165:14]
  assign _GEN_21 = _T_56 ? output_ : 32'h0; // @[Conditional.scala 39:67]
  assign _GEN_30 = _T_52 ? 1'h0 : _T_56; // @[Conditional.scala 39:67]
  assign _GEN_32 = _T_52 ? 32'h0 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_50 ? _GEN_8 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_41 = _T_50 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_43 = _T_50 ? 32'h0 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_48 = _T_48 ? _GEN_6 : _GEN_36; // @[Conditional.scala 40:58]
  assign io_NodeReq_ready = state == 2'h0; // @[ReadMemoryController.scala 83:20]
  assign io_MemReq_valid = _T_48 ? 1'h0 : _T_50; // @[ReadMemoryController.scala 95:19 ReadMemoryController.scala 140:23]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_57; // @[ReadMemoryController.scala 96:23]
  assign io_MemReq_bits_tag = {{7'd0}, ID}; // @[ReadMemoryController.scala 99:22]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[ReadMemoryController.scala 104:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[ReadMemoryController.scala 101:26]
  assign io_output_valid = _T_48 ? 1'h0 : _GEN_41; // @[ReadMemoryController.scala 90:19 ReadMemoryController.scala 164:23]
  assign io_output_bits_RouteID = request_R_RouteID; // @[ReadMemoryController.scala 91:26]
  assign io_output_bits_data = _T_48 ? 32'h0 : _GEN_43; // @[ReadMemoryController.scala 93:23 ReadMemoryController.scala 168:29]
  assign io_free = state == 2'h0; // @[ReadMemoryController.scala 81:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ID = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_RouteID = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  request_R_address = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  request_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {2{`RANDOM}};
  bitmask = _RAND_4[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  sendbytemask = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ReqAddress = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ptr = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  linebuffer_0 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  linebuffer_1 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  isWrite = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      ID <= 1'h0;
    end else begin
      ID <= 1'h1;
    end
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_9) begin
        request_R_RouteID <= io_NodeReq_bits_RouteID;
      end
    end
    if (reset) begin
      request_R_address <= 32'h0;
    end else begin
      if (_T_9) begin
        request_R_address <= io_NodeReq_bits_address;
      end
    end
    if (reset) begin
      request_R_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      bitmask <= 64'h0;
    end else begin
      bitmask <= _GEN_5[63:0];
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_48[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_9) begin
        ReqAddress <= _T_11;
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              ptr <= _T_54;
            end
          end else begin
            if (_T_56) begin
              ptr <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (1'h0 == ptr) begin
                linebuffer_0 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (ptr) begin
                linebuffer_1 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_48) begin
        if (_T_9) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_50) begin
          if (io_MemReq_ready) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (_T_55) begin
                state <= 2'h3;
              end else begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_56) begin
              if (io_output_ready) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    isWrite <= reset;
  end
endmodule
module ReadMemoryController(
  input         clock,
  input         reset,
  output        io_ReadIn_0_ready,
  input         io_ReadIn_0_valid,
  input  [31:0] io_ReadIn_0_bits_address,
  input  [4:0]  io_ReadIn_0_bits_taskID,
  output        io_ReadIn_1_ready,
  input         io_ReadIn_1_valid,
  input  [31:0] io_ReadIn_1_bits_address,
  input  [4:0]  io_ReadIn_1_bits_taskID,
  output        io_ReadOut_0_valid,
  output [31:0] io_ReadOut_0_data,
  output        io_ReadOut_1_valid,
  output [31:0] io_ReadOut_1_data,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag
);
  wire  in_arb_clock; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_0_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_0_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_0_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_0_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_1_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_1_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_1_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_1_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_out_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_out_valid; // @[ReadMemoryController.scala 221:25]
  wire [15:0] in_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_out_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  alloc_arb_io_in_0_ready; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_in_0_valid; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_in_1_ready; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_in_1_valid; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_out_ready; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_out_valid; // @[ReadMemoryController.scala 223:25]
  wire  cachereq_arb_io_in_0_ready; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_0_valid; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_0_bits_addr; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_0_bits_data; // @[ReadMemoryController.scala 226:31]
  wire [3:0] cachereq_arb_io_in_0_bits_mask; // @[ReadMemoryController.scala 226:31]
  wire [7:0] cachereq_arb_io_in_0_bits_tag; // @[ReadMemoryController.scala 226:31]
  wire [4:0] cachereq_arb_io_in_0_bits_taskID; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_0_bits_iswrite; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_1_ready; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_1_valid; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_1_bits_addr; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_1_bits_data; // @[ReadMemoryController.scala 226:31]
  wire [3:0] cachereq_arb_io_in_1_bits_mask; // @[ReadMemoryController.scala 226:31]
  wire [7:0] cachereq_arb_io_in_1_bits_tag; // @[ReadMemoryController.scala 226:31]
  wire [4:0] cachereq_arb_io_in_1_bits_taskID; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_1_bits_iswrite; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_out_ready; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_out_valid; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_out_bits_addr; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_out_bits_data; // @[ReadMemoryController.scala 226:31]
  wire [3:0] cachereq_arb_io_out_bits_mask; // @[ReadMemoryController.scala 226:31]
  wire [7:0] cachereq_arb_io_out_bits_tag; // @[ReadMemoryController.scala 226:31]
  wire [4:0] cachereq_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_out_bits_iswrite; // @[ReadMemoryController.scala 226:31]
  wire  cacheresp_demux_io_en; // @[ReadMemoryController.scala 228:31]
  wire [31:0] cacheresp_demux_io_input_data; // @[ReadMemoryController.scala 228:31]
  wire [7:0] cacheresp_demux_io_input_tag; // @[ReadMemoryController.scala 228:31]
  wire  cacheresp_demux_io_sel; // @[ReadMemoryController.scala 228:31]
  wire  cacheresp_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 228:31]
  wire [31:0] cacheresp_demux_io_outputs_0_data; // @[ReadMemoryController.scala 228:31]
  wire [7:0] cacheresp_demux_io_outputs_0_tag; // @[ReadMemoryController.scala 228:31]
  wire  cacheresp_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 228:31]
  wire [31:0] cacheresp_demux_io_outputs_1_data; // @[ReadMemoryController.scala 228:31]
  wire [7:0] cacheresp_demux_io_outputs_1_tag; // @[ReadMemoryController.scala 228:31]
  wire  out_arb_clock; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_0_ready; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_0_valid; // @[ReadMemoryController.scala 231:25]
  wire [15:0] out_arb_io_in_0_bits_RouteID; // @[ReadMemoryController.scala 231:25]
  wire [31:0] out_arb_io_in_0_bits_data; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_1_ready; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_1_valid; // @[ReadMemoryController.scala 231:25]
  wire [15:0] out_arb_io_in_1_bits_RouteID; // @[ReadMemoryController.scala 231:25]
  wire [31:0] out_arb_io_in_1_bits_data; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_out_ready; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_out_valid; // @[ReadMemoryController.scala 231:25]
  wire [15:0] out_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 231:25]
  wire [31:0] out_arb_io_out_bits_data; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_chosen; // @[ReadMemoryController.scala 231:25]
  wire  out_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_0_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_1_data; // @[ReadMemoryController.scala 232:25]
  wire [15:0] out_demux_io_input_RouteID; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_input_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_enable; // @[ReadMemoryController.scala 232:25]
  wire  ReadTable_0_clock; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_reset; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_NodeReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_NodeReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_0_io_NodeReq_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_NodeReq_bits_address; // @[ReadMemoryController.scala 251:28]
  wire [4:0] ReadTable_0_io_NodeReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_MemReq_bits_addr; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_0_io_MemReq_bits_tag; // @[ReadMemoryController.scala 251:28]
  wire [4:0] ReadTable_0_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemResp_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_MemResp_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_output_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_output_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_0_io_output_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_output_bits_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_free; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_clock; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_reset; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_NodeReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_NodeReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_1_io_NodeReq_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_NodeReq_bits_address; // @[ReadMemoryController.scala 251:28]
  wire [4:0] ReadTable_1_io_NodeReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_MemReq_bits_addr; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_1_io_MemReq_bits_tag; // @[ReadMemoryController.scala 251:28]
  wire [4:0] ReadTable_1_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemResp_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_MemResp_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_output_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_output_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_1_io_output_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_output_bits_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_free; // @[ReadMemoryController.scala 251:28]
  ArbiterTree_1 in_arb ( // @[ReadMemoryController.scala 221:25]
    .clock(in_arb_clock),
    .io_in_0_ready(in_arb_io_in_0_ready),
    .io_in_0_valid(in_arb_io_in_0_valid),
    .io_in_0_bits_address(in_arb_io_in_0_bits_address),
    .io_in_0_bits_taskID(in_arb_io_in_0_bits_taskID),
    .io_in_1_ready(in_arb_io_in_1_ready),
    .io_in_1_valid(in_arb_io_in_1_valid),
    .io_in_1_bits_address(in_arb_io_in_1_bits_address),
    .io_in_1_bits_taskID(in_arb_io_in_1_bits_taskID),
    .io_out_ready(in_arb_io_out_ready),
    .io_out_valid(in_arb_io_out_valid),
    .io_out_bits_RouteID(in_arb_io_out_bits_RouteID),
    .io_out_bits_address(in_arb_io_out_bits_address),
    .io_out_bits_taskID(in_arb_io_out_bits_taskID)
  );
  Arbiter alloc_arb ( // @[ReadMemoryController.scala 223:25]
    .io_in_0_ready(alloc_arb_io_in_0_ready),
    .io_in_0_valid(alloc_arb_io_in_0_valid),
    .io_in_1_ready(alloc_arb_io_in_1_ready),
    .io_in_1_valid(alloc_arb_io_in_1_valid),
    .io_out_ready(alloc_arb_io_out_ready),
    .io_out_valid(alloc_arb_io_out_valid)
  );
  Arbiter_1 cachereq_arb ( // @[ReadMemoryController.scala 226:31]
    .io_in_0_ready(cachereq_arb_io_in_0_ready),
    .io_in_0_valid(cachereq_arb_io_in_0_valid),
    .io_in_0_bits_addr(cachereq_arb_io_in_0_bits_addr),
    .io_in_0_bits_data(cachereq_arb_io_in_0_bits_data),
    .io_in_0_bits_mask(cachereq_arb_io_in_0_bits_mask),
    .io_in_0_bits_tag(cachereq_arb_io_in_0_bits_tag),
    .io_in_0_bits_taskID(cachereq_arb_io_in_0_bits_taskID),
    .io_in_0_bits_iswrite(cachereq_arb_io_in_0_bits_iswrite),
    .io_in_1_ready(cachereq_arb_io_in_1_ready),
    .io_in_1_valid(cachereq_arb_io_in_1_valid),
    .io_in_1_bits_addr(cachereq_arb_io_in_1_bits_addr),
    .io_in_1_bits_data(cachereq_arb_io_in_1_bits_data),
    .io_in_1_bits_mask(cachereq_arb_io_in_1_bits_mask),
    .io_in_1_bits_tag(cachereq_arb_io_in_1_bits_tag),
    .io_in_1_bits_taskID(cachereq_arb_io_in_1_bits_taskID),
    .io_in_1_bits_iswrite(cachereq_arb_io_in_1_bits_iswrite),
    .io_out_ready(cachereq_arb_io_out_ready),
    .io_out_valid(cachereq_arb_io_out_valid),
    .io_out_bits_addr(cachereq_arb_io_out_bits_addr),
    .io_out_bits_data(cachereq_arb_io_out_bits_data),
    .io_out_bits_mask(cachereq_arb_io_out_bits_mask),
    .io_out_bits_tag(cachereq_arb_io_out_bits_tag),
    .io_out_bits_taskID(cachereq_arb_io_out_bits_taskID),
    .io_out_bits_iswrite(cachereq_arb_io_out_bits_iswrite)
  );
  Demux cacheresp_demux ( // @[ReadMemoryController.scala 228:31]
    .io_en(cacheresp_demux_io_en),
    .io_input_data(cacheresp_demux_io_input_data),
    .io_input_tag(cacheresp_demux_io_input_tag),
    .io_sel(cacheresp_demux_io_sel),
    .io_outputs_0_valid(cacheresp_demux_io_outputs_0_valid),
    .io_outputs_0_data(cacheresp_demux_io_outputs_0_data),
    .io_outputs_0_tag(cacheresp_demux_io_outputs_0_tag),
    .io_outputs_1_valid(cacheresp_demux_io_outputs_1_valid),
    .io_outputs_1_data(cacheresp_demux_io_outputs_1_data),
    .io_outputs_1_tag(cacheresp_demux_io_outputs_1_tag)
  );
  RRArbiter_1 out_arb ( // @[ReadMemoryController.scala 231:25]
    .clock(out_arb_clock),
    .io_in_0_ready(out_arb_io_in_0_ready),
    .io_in_0_valid(out_arb_io_in_0_valid),
    .io_in_0_bits_RouteID(out_arb_io_in_0_bits_RouteID),
    .io_in_0_bits_data(out_arb_io_in_0_bits_data),
    .io_in_1_ready(out_arb_io_in_1_ready),
    .io_in_1_valid(out_arb_io_in_1_valid),
    .io_in_1_bits_RouteID(out_arb_io_in_1_bits_RouteID),
    .io_in_1_bits_data(out_arb_io_in_1_bits_data),
    .io_out_ready(out_arb_io_out_ready),
    .io_out_valid(out_arb_io_out_valid),
    .io_out_bits_RouteID(out_arb_io_out_bits_RouteID),
    .io_out_bits_data(out_arb_io_out_bits_data),
    .io_chosen(out_arb_io_chosen)
  );
  DeMuxTree_1 out_demux ( // @[ReadMemoryController.scala 232:25]
    .io_outputs_0_valid(out_demux_io_outputs_0_valid),
    .io_outputs_0_data(out_demux_io_outputs_0_data),
    .io_outputs_1_valid(out_demux_io_outputs_1_valid),
    .io_outputs_1_data(out_demux_io_outputs_1_data),
    .io_input_RouteID(out_demux_io_input_RouteID),
    .io_input_data(out_demux_io_input_data),
    .io_enable(out_demux_io_enable)
  );
  ReadTableEntry ReadTable_0 ( // @[ReadMemoryController.scala 251:28]
    .clock(ReadTable_0_clock),
    .reset(ReadTable_0_reset),
    .io_NodeReq_ready(ReadTable_0_io_NodeReq_ready),
    .io_NodeReq_valid(ReadTable_0_io_NodeReq_valid),
    .io_NodeReq_bits_RouteID(ReadTable_0_io_NodeReq_bits_RouteID),
    .io_NodeReq_bits_address(ReadTable_0_io_NodeReq_bits_address),
    .io_NodeReq_bits_taskID(ReadTable_0_io_NodeReq_bits_taskID),
    .io_MemReq_ready(ReadTable_0_io_MemReq_ready),
    .io_MemReq_valid(ReadTable_0_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadTable_0_io_MemReq_bits_addr),
    .io_MemReq_bits_tag(ReadTable_0_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadTable_0_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadTable_0_io_MemReq_bits_iswrite),
    .io_MemResp_valid(ReadTable_0_io_MemResp_valid),
    .io_MemResp_data(ReadTable_0_io_MemResp_data),
    .io_output_ready(ReadTable_0_io_output_ready),
    .io_output_valid(ReadTable_0_io_output_valid),
    .io_output_bits_RouteID(ReadTable_0_io_output_bits_RouteID),
    .io_output_bits_data(ReadTable_0_io_output_bits_data),
    .io_free(ReadTable_0_io_free)
  );
  ReadTableEntry_1 ReadTable_1 ( // @[ReadMemoryController.scala 251:28]
    .clock(ReadTable_1_clock),
    .reset(ReadTable_1_reset),
    .io_NodeReq_ready(ReadTable_1_io_NodeReq_ready),
    .io_NodeReq_valid(ReadTable_1_io_NodeReq_valid),
    .io_NodeReq_bits_RouteID(ReadTable_1_io_NodeReq_bits_RouteID),
    .io_NodeReq_bits_address(ReadTable_1_io_NodeReq_bits_address),
    .io_NodeReq_bits_taskID(ReadTable_1_io_NodeReq_bits_taskID),
    .io_MemReq_ready(ReadTable_1_io_MemReq_ready),
    .io_MemReq_valid(ReadTable_1_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadTable_1_io_MemReq_bits_addr),
    .io_MemReq_bits_tag(ReadTable_1_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadTable_1_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadTable_1_io_MemReq_bits_iswrite),
    .io_MemResp_valid(ReadTable_1_io_MemResp_valid),
    .io_MemResp_data(ReadTable_1_io_MemResp_data),
    .io_output_ready(ReadTable_1_io_output_ready),
    .io_output_valid(ReadTable_1_io_output_valid),
    .io_output_bits_RouteID(ReadTable_1_io_output_bits_RouteID),
    .io_output_bits_data(ReadTable_1_io_output_bits_data),
    .io_free(ReadTable_1_io_free)
  );
  assign io_ReadIn_0_ready = in_arb_io_in_0_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_1_ready = in_arb_io_in_1_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadOut_0_valid = out_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_0_data = out_demux_io_outputs_0_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_1_valid = out_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_1_data = out_demux_io_outputs_1_data; // @[ReadMemoryController.scala 241:19]
  assign io_MemReq_valid = cachereq_arb_io_out_valid; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_addr = cachereq_arb_io_out_bits_addr; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_data = cachereq_arb_io_out_bits_data; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_mask = cachereq_arb_io_out_bits_mask; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_tag = cachereq_arb_io_out_bits_tag; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_taskID = cachereq_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_iswrite = cachereq_arb_io_out_bits_iswrite; // @[ReadMemoryController.scala 288:13]
  assign in_arb_clock = clock;
  assign in_arb_io_in_0_valid = io_ReadIn_0_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_0_bits_address = io_ReadIn_0_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_0_bits_taskID = io_ReadIn_0_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_1_valid = io_ReadIn_1_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_1_bits_address = io_ReadIn_1_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_1_bits_taskID = io_ReadIn_1_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_out_ready = alloc_arb_io_out_valid; // @[ReadMemoryController.scala 283:23]
  assign alloc_arb_io_in_0_valid = ReadTable_0_io_free; // @[ReadMemoryController.scala 254:30]
  assign alloc_arb_io_in_1_valid = ReadTable_1_io_free; // @[ReadMemoryController.scala 254:30]
  assign alloc_arb_io_out_ready = in_arb_io_out_valid; // @[ReadMemoryController.scala 284:26]
  assign cachereq_arb_io_in_0_valid = ReadTable_0_io_MemReq_valid; // @[ReadMemoryController.scala 260:33]
  assign cachereq_arb_io_in_0_bits_addr = ReadTable_0_io_MemReq_bits_addr; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_data = 32'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_mask = 4'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_tag = ReadTable_0_io_MemReq_bits_tag; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_taskID = ReadTable_0_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_iswrite = ReadTable_0_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_valid = ReadTable_1_io_MemReq_valid; // @[ReadMemoryController.scala 260:33]
  assign cachereq_arb_io_in_1_bits_addr = ReadTable_1_io_MemReq_bits_addr; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_data = 32'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_mask = 4'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_tag = ReadTable_1_io_MemReq_bits_tag; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_taskID = ReadTable_1_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_iswrite = ReadTable_1_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_out_ready = io_MemReq_ready; // @[ReadMemoryController.scala 288:13]
  assign cacheresp_demux_io_en = io_MemResp_valid; // @[ReadMemoryController.scala 291:25]
  assign cacheresp_demux_io_input_data = io_MemResp_bits_data; // @[ReadMemoryController.scala 292:28]
  assign cacheresp_demux_io_input_tag = io_MemResp_bits_tag; // @[ReadMemoryController.scala 292:28]
  assign cacheresp_demux_io_sel = io_MemResp_bits_tag[0]; // @[ReadMemoryController.scala 293:26]
  assign out_arb_clock = clock;
  assign out_arb_io_in_0_valid = ReadTable_0_io_output_valid; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_0_bits_RouteID = ReadTable_0_io_output_bits_RouteID; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_0_bits_data = ReadTable_0_io_output_bits_data; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_1_valid = ReadTable_1_io_output_valid; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_1_bits_RouteID = ReadTable_1_io_output_bits_RouteID; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_1_bits_data = ReadTable_1_io_output_bits_data; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_out_ready = 1'h1; // @[ReadMemoryController.scala 296:24]
  assign out_demux_io_input_RouteID = out_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 298:22]
  assign out_demux_io_input_data = out_arb_io_out_bits_data; // @[ReadMemoryController.scala 298:22]
  assign out_demux_io_enable = out_arb_io_out_ready & out_arb_io_out_valid; // @[ReadMemoryController.scala 297:23]
  assign ReadTable_0_clock = clock;
  assign ReadTable_0_reset = reset;
  assign ReadTable_0_io_NodeReq_valid = alloc_arb_io_in_0_ready & alloc_arb_io_in_0_valid; // @[ReadMemoryController.scala 256:33]
  assign ReadTable_0_io_NodeReq_bits_RouteID = in_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_MemReq_ready = cachereq_arb_io_in_0_ready; // @[ReadMemoryController.scala 262:32]
  assign ReadTable_0_io_MemResp_valid = cacheresp_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_0_io_MemResp_data = cacheresp_demux_io_outputs_0_data; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_0_io_output_ready = out_arb_io_in_0_ready; // @[ReadMemoryController.scala 268:22]
  assign ReadTable_1_clock = clock;
  assign ReadTable_1_reset = reset;
  assign ReadTable_1_io_NodeReq_valid = alloc_arb_io_in_1_ready & alloc_arb_io_in_1_valid; // @[ReadMemoryController.scala 256:33]
  assign ReadTable_1_io_NodeReq_bits_RouteID = in_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_MemReq_ready = cachereq_arb_io_in_1_ready; // @[ReadMemoryController.scala 262:32]
  assign ReadTable_1_io_MemResp_valid = cacheresp_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_1_io_MemResp_data = cacheresp_demux_io_outputs_1_data; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_1_io_output_ready = out_arb_io_in_1_ready; // @[ReadMemoryController.scala 268:22]
endmodule
module RRArbiter_2(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [31:0] io_in_0_bits_data,
  input  [3:0]  io_in_0_bits_mask,
  input  [7:0]  io_in_0_bits_tag,
  input  [4:0]  io_in_0_bits_taskID,
  input         io_in_0_bits_iswrite,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [31:0] io_in_1_bits_data,
  input  [3:0]  io_in_1_bits_mask,
  input  [7:0]  io_in_1_bits_tag,
  input  [4:0]  io_in_1_bits_taskID,
  input         io_in_1_bits_iswrite,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [31:0] io_out_bits_data,
  output [3:0]  io_out_bits_mask,
  output [7:0]  io_out_bits_tag,
  output [4:0]  io_out_bits_taskID,
  output        io_out_bits_iswrite,
  output        io_chosen
);
  wire  _T; // @[Decoupled.scala 40:37]
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Arbiter.scala 67:57]
  wire  _T_5; // @[Arbiter.scala 68:83]
  wire  _T_7; // @[Arbiter.scala 31:68]
  wire  _T_9; // @[Arbiter.scala 31:78]
  wire  _T_10; // @[Arbiter.scala 31:78]
  wire  _T_14; // @[Arbiter.scala 72:50]
  wire  _GEN_19; // @[Arbiter.scala 77:27]
  assign _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = 1'h1 > _T_1; // @[Arbiter.scala 67:57]
  assign _T_5 = io_in_1_valid & _T_3; // @[Arbiter.scala 68:83]
  assign _T_7 = _T_5 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_9 = _T_5 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_10 = _T_7 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_14 = _T_3 | _T_10; // @[Arbiter.scala 72:50]
  assign _GEN_19 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_9 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_14 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_out_bits_mask = io_chosen ? io_in_1_bits_mask : io_in_0_bits_mask; // @[Arbiter.scala 42:15]
  assign io_out_bits_tag = io_chosen ? io_in_1_bits_tag : io_in_0_bits_tag; // @[Arbiter.scala 42:15]
  assign io_out_bits_taskID = io_chosen ? io_in_1_bits_taskID : io_in_0_bits_taskID; // @[Arbiter.scala 42:15]
  assign io_out_bits_iswrite = io_chosen ? io_in_1_bits_iswrite : io_in_0_bits_iswrite; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_5 | _GEN_19; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (_T) begin
      _T_1 <= io_chosen;
    end
  end
endmodule
module ReadWriteArbiter(
  input         clock,
  output        io_ReadMemReq_ready,
  input         io_ReadMemReq_valid,
  input  [31:0] io_ReadMemReq_bits_addr,
  input  [31:0] io_ReadMemReq_bits_data,
  input  [3:0]  io_ReadMemReq_bits_mask,
  input  [7:0]  io_ReadMemReq_bits_tag,
  input  [4:0]  io_ReadMemReq_bits_taskID,
  input         io_ReadMemReq_bits_iswrite,
  output        io_WriteMemReq_ready,
  input         io_WriteMemReq_valid,
  input  [31:0] io_WriteMemReq_bits_addr,
  input  [31:0] io_WriteMemReq_bits_data,
  input  [3:0]  io_WriteMemReq_bits_mask,
  input  [7:0]  io_WriteMemReq_bits_tag,
  input  [4:0]  io_WriteMemReq_bits_taskID,
  input         io_WriteMemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemResp_bits_iswrite,
  output        io_ReadMemResp_valid,
  output [31:0] io_ReadMemResp_bits_data,
  output [7:0]  io_ReadMemResp_bits_tag,
  output        io_WriteMemResp_valid,
  output [31:0] io_WriteMemResp_bits_data,
  output [7:0]  io_WriteMemResp_bits_tag,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite
);
  wire  cachereq_arb_clock; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_0_ready; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_0_valid; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_0_bits_addr; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_0_bits_data; // @[ReadWriteArbiter.scala 48:31]
  wire [3:0] cachereq_arb_io_in_0_bits_mask; // @[ReadWriteArbiter.scala 48:31]
  wire [7:0] cachereq_arb_io_in_0_bits_tag; // @[ReadWriteArbiter.scala 48:31]
  wire [4:0] cachereq_arb_io_in_0_bits_taskID; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_0_bits_iswrite; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_1_ready; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_1_valid; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_1_bits_addr; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_1_bits_data; // @[ReadWriteArbiter.scala 48:31]
  wire [3:0] cachereq_arb_io_in_1_bits_mask; // @[ReadWriteArbiter.scala 48:31]
  wire [7:0] cachereq_arb_io_in_1_bits_tag; // @[ReadWriteArbiter.scala 48:31]
  wire [4:0] cachereq_arb_io_in_1_bits_taskID; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_1_bits_iswrite; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_out_ready; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_out_valid; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_out_bits_addr; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_out_bits_data; // @[ReadWriteArbiter.scala 48:31]
  wire [3:0] cachereq_arb_io_out_bits_mask; // @[ReadWriteArbiter.scala 48:31]
  wire [7:0] cachereq_arb_io_out_bits_tag; // @[ReadWriteArbiter.scala 48:31]
  wire [4:0] cachereq_arb_io_out_bits_taskID; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_out_bits_iswrite; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_chosen; // @[ReadWriteArbiter.scala 48:31]
  wire  cacheresp_demux_io_en; // @[ReadWriteArbiter.scala 50:31]
  wire [31:0] cacheresp_demux_io_input_data; // @[ReadWriteArbiter.scala 50:31]
  wire [7:0] cacheresp_demux_io_input_tag; // @[ReadWriteArbiter.scala 50:31]
  wire  cacheresp_demux_io_sel; // @[ReadWriteArbiter.scala 50:31]
  wire  cacheresp_demux_io_outputs_0_valid; // @[ReadWriteArbiter.scala 50:31]
  wire [31:0] cacheresp_demux_io_outputs_0_data; // @[ReadWriteArbiter.scala 50:31]
  wire [7:0] cacheresp_demux_io_outputs_0_tag; // @[ReadWriteArbiter.scala 50:31]
  wire  cacheresp_demux_io_outputs_1_valid; // @[ReadWriteArbiter.scala 50:31]
  wire [31:0] cacheresp_demux_io_outputs_1_data; // @[ReadWriteArbiter.scala 50:31]
  wire [7:0] cacheresp_demux_io_outputs_1_tag; // @[ReadWriteArbiter.scala 50:31]
  RRArbiter_2 cachereq_arb ( // @[ReadWriteArbiter.scala 48:31]
    .clock(cachereq_arb_clock),
    .io_in_0_ready(cachereq_arb_io_in_0_ready),
    .io_in_0_valid(cachereq_arb_io_in_0_valid),
    .io_in_0_bits_addr(cachereq_arb_io_in_0_bits_addr),
    .io_in_0_bits_data(cachereq_arb_io_in_0_bits_data),
    .io_in_0_bits_mask(cachereq_arb_io_in_0_bits_mask),
    .io_in_0_bits_tag(cachereq_arb_io_in_0_bits_tag),
    .io_in_0_bits_taskID(cachereq_arb_io_in_0_bits_taskID),
    .io_in_0_bits_iswrite(cachereq_arb_io_in_0_bits_iswrite),
    .io_in_1_ready(cachereq_arb_io_in_1_ready),
    .io_in_1_valid(cachereq_arb_io_in_1_valid),
    .io_in_1_bits_addr(cachereq_arb_io_in_1_bits_addr),
    .io_in_1_bits_data(cachereq_arb_io_in_1_bits_data),
    .io_in_1_bits_mask(cachereq_arb_io_in_1_bits_mask),
    .io_in_1_bits_tag(cachereq_arb_io_in_1_bits_tag),
    .io_in_1_bits_taskID(cachereq_arb_io_in_1_bits_taskID),
    .io_in_1_bits_iswrite(cachereq_arb_io_in_1_bits_iswrite),
    .io_out_ready(cachereq_arb_io_out_ready),
    .io_out_valid(cachereq_arb_io_out_valid),
    .io_out_bits_addr(cachereq_arb_io_out_bits_addr),
    .io_out_bits_data(cachereq_arb_io_out_bits_data),
    .io_out_bits_mask(cachereq_arb_io_out_bits_mask),
    .io_out_bits_tag(cachereq_arb_io_out_bits_tag),
    .io_out_bits_taskID(cachereq_arb_io_out_bits_taskID),
    .io_out_bits_iswrite(cachereq_arb_io_out_bits_iswrite),
    .io_chosen(cachereq_arb_io_chosen)
  );
  Demux cacheresp_demux ( // @[ReadWriteArbiter.scala 50:31]
    .io_en(cacheresp_demux_io_en),
    .io_input_data(cacheresp_demux_io_input_data),
    .io_input_tag(cacheresp_demux_io_input_tag),
    .io_sel(cacheresp_demux_io_sel),
    .io_outputs_0_valid(cacheresp_demux_io_outputs_0_valid),
    .io_outputs_0_data(cacheresp_demux_io_outputs_0_data),
    .io_outputs_0_tag(cacheresp_demux_io_outputs_0_tag),
    .io_outputs_1_valid(cacheresp_demux_io_outputs_1_valid),
    .io_outputs_1_data(cacheresp_demux_io_outputs_1_data),
    .io_outputs_1_tag(cacheresp_demux_io_outputs_1_tag)
  );
  assign io_ReadMemReq_ready = cachereq_arb_io_in_0_ready; // @[ReadWriteArbiter.scala 57:29]
  assign io_WriteMemReq_ready = cachereq_arb_io_in_1_ready; // @[ReadWriteArbiter.scala 58:29]
  assign io_ReadMemResp_valid = cacheresp_demux_io_outputs_0_valid; // @[ReadWriteArbiter.scala 69:24]
  assign io_ReadMemResp_bits_data = cacheresp_demux_io_outputs_0_data; // @[ReadWriteArbiter.scala 68:23]
  assign io_ReadMemResp_bits_tag = cacheresp_demux_io_outputs_0_tag; // @[ReadWriteArbiter.scala 68:23]
  assign io_WriteMemResp_valid = cacheresp_demux_io_outputs_1_valid; // @[ReadWriteArbiter.scala 71:25]
  assign io_WriteMemResp_bits_data = cacheresp_demux_io_outputs_1_data; // @[ReadWriteArbiter.scala 70:24]
  assign io_WriteMemResp_bits_tag = cacheresp_demux_io_outputs_1_tag; // @[ReadWriteArbiter.scala 70:24]
  assign io_MemReq_valid = cachereq_arb_io_out_valid; // @[ReadWriteArbiter.scala 62:19]
  assign io_MemReq_bits_addr = cachereq_arb_io_out_bits_addr; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_data = cachereq_arb_io_out_bits_data; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_mask = cachereq_arb_io_out_bits_mask; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_tag = cachereq_arb_io_out_bits_tag; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_taskID = cachereq_arb_io_out_bits_taskID; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_iswrite = cachereq_arb_io_out_bits_iswrite; // @[ReadWriteArbiter.scala 61:18]
  assign cachereq_arb_clock = clock;
  assign cachereq_arb_io_in_0_valid = io_ReadMemReq_valid; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_addr = io_ReadMemReq_bits_addr; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_data = io_ReadMemReq_bits_data; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_mask = io_ReadMemReq_bits_mask; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_tag = io_ReadMemReq_bits_tag; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_taskID = io_ReadMemReq_bits_taskID; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_iswrite = io_ReadMemReq_bits_iswrite; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_1_valid = io_WriteMemReq_valid; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_addr = io_WriteMemReq_bits_addr; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_data = io_WriteMemReq_bits_data; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_mask = io_WriteMemReq_bits_mask; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_tag = io_WriteMemReq_bits_tag; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_taskID = io_WriteMemReq_bits_taskID; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_iswrite = io_WriteMemReq_bits_iswrite; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_out_ready = io_MemReq_ready; // @[ReadWriteArbiter.scala 60:29]
  assign cacheresp_demux_io_en = io_MemResp_valid; // @[ReadWriteArbiter.scala 76:25]
  assign cacheresp_demux_io_input_data = io_MemResp_bits_data; // @[ReadWriteArbiter.scala 77:28]
  assign cacheresp_demux_io_input_tag = io_MemResp_bits_tag; // @[ReadWriteArbiter.scala 77:28]
  assign cacheresp_demux_io_sel = io_MemResp_bits_iswrite; // @[ReadWriteArbiter.scala 80:26]
endmodule
module UnifiedController(
  input         clock,
  input         reset,
  output        io_WriteIn_0_ready,
  input         io_WriteIn_0_valid,
  input  [21:0] io_WriteIn_0_bits_address,
  input  [31:0] io_WriteIn_0_bits_data,
  input  [4:0]  io_WriteIn_0_bits_taskID,
  output        io_WriteOut_0_valid,
  output        io_ReadIn_0_ready,
  input         io_ReadIn_0_valid,
  input  [31:0] io_ReadIn_0_bits_address,
  input  [4:0]  io_ReadIn_0_bits_taskID,
  output        io_ReadIn_1_ready,
  input         io_ReadIn_1_valid,
  input  [31:0] io_ReadIn_1_bits_address,
  input  [4:0]  io_ReadIn_1_bits_taskID,
  output        io_ReadOut_0_valid,
  output [31:0] io_ReadOut_0_data,
  output        io_ReadOut_1_valid,
  output [31:0] io_ReadOut_1_data,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemResp_bits_iswrite,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite
);
  wire  WriteController_clock; // @[UnifiedController.scala 53:32]
  wire  WriteController_reset; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_0_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_0_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_0_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_0_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_0_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_0_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_MemReq_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_MemReq_valid; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_MemReq_bits_addr; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_MemReq_bits_data; // @[UnifiedController.scala 53:32]
  wire [3:0] WriteController_io_MemReq_bits_mask; // @[UnifiedController.scala 53:32]
  wire [7:0] WriteController_io_MemReq_bits_tag; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_MemReq_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_MemResp_valid; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_MemResp_bits_data; // @[UnifiedController.scala 53:32]
  wire [7:0] WriteController_io_MemResp_bits_tag; // @[UnifiedController.scala 53:32]
  wire  ReadController_clock; // @[UnifiedController.scala 54:32]
  wire  ReadController_reset; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_0_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_0_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_0_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_0_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_1_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_1_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_1_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_1_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_0_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_0_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_1_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_1_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_MemReq_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_MemReq_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_MemReq_bits_addr; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_MemReq_bits_data; // @[UnifiedController.scala 54:32]
  wire [3:0] ReadController_io_MemReq_bits_mask; // @[UnifiedController.scala 54:32]
  wire [7:0] ReadController_io_MemReq_bits_tag; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_MemReq_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_MemResp_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_MemResp_bits_data; // @[UnifiedController.scala 54:32]
  wire [7:0] ReadController_io_MemResp_bits_tag; // @[UnifiedController.scala 54:32]
  wire  ReadWriteArbiter_clock; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_ReadMemReq_ready; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_ReadMemReq_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_ReadMemReq_bits_addr; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_ReadMemReq_bits_data; // @[UnifiedController.scala 55:32]
  wire [3:0] ReadWriteArbiter_io_ReadMemReq_bits_mask; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_ReadMemReq_bits_tag; // @[UnifiedController.scala 55:32]
  wire [4:0] ReadWriteArbiter_io_ReadMemReq_bits_taskID; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_ReadMemReq_bits_iswrite; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_WriteMemReq_ready; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_WriteMemReq_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_WriteMemReq_bits_addr; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_WriteMemReq_bits_data; // @[UnifiedController.scala 55:32]
  wire [3:0] ReadWriteArbiter_io_WriteMemReq_bits_mask; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_WriteMemReq_bits_tag; // @[UnifiedController.scala 55:32]
  wire [4:0] ReadWriteArbiter_io_WriteMemReq_bits_taskID; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_WriteMemReq_bits_iswrite; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemResp_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_MemResp_bits_data; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_MemResp_bits_tag; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemResp_bits_iswrite; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_ReadMemResp_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_ReadMemResp_bits_data; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_ReadMemResp_bits_tag; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_WriteMemResp_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_WriteMemResp_bits_data; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_WriteMemResp_bits_tag; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemReq_ready; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemReq_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_MemReq_bits_addr; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_MemReq_bits_data; // @[UnifiedController.scala 55:32]
  wire [3:0] ReadWriteArbiter_io_MemReq_bits_mask; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_MemReq_bits_tag; // @[UnifiedController.scala 55:32]
  wire [4:0] ReadWriteArbiter_io_MemReq_bits_taskID; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemReq_bits_iswrite; // @[UnifiedController.scala 55:32]
  wire  _T; // @[Decoupled.scala 40:37]
  wire  _T_1; // @[UnifiedController.scala 92:15]
  wire  _T_2; // @[UnifiedController.scala 92:15]
  wire  _GEN_0; // @[UnifiedController.scala 92:15]
  wire  _GEN_1; // @[UnifiedController.scala 94:15]
  wire  _GEN_2; // @[UnifiedController.scala 94:15]
  wire  _GEN_3; // @[UnifiedController.scala 100:15]
  wire  _GEN_4; // @[UnifiedController.scala 102:15]
  wire  _GEN_5; // @[UnifiedController.scala 102:15]
  WriteMemoryController WriteController ( // @[UnifiedController.scala 53:32]
    .clock(WriteController_clock),
    .reset(WriteController_reset),
    .io_WriteIn_0_ready(WriteController_io_WriteIn_0_ready),
    .io_WriteIn_0_valid(WriteController_io_WriteIn_0_valid),
    .io_WriteIn_0_bits_address(WriteController_io_WriteIn_0_bits_address),
    .io_WriteIn_0_bits_data(WriteController_io_WriteIn_0_bits_data),
    .io_WriteIn_0_bits_taskID(WriteController_io_WriteIn_0_bits_taskID),
    .io_WriteOut_0_valid(WriteController_io_WriteOut_0_valid),
    .io_MemReq_ready(WriteController_io_MemReq_ready),
    .io_MemReq_valid(WriteController_io_MemReq_valid),
    .io_MemReq_bits_addr(WriteController_io_MemReq_bits_addr),
    .io_MemReq_bits_data(WriteController_io_MemReq_bits_data),
    .io_MemReq_bits_mask(WriteController_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(WriteController_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(WriteController_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(WriteController_io_MemReq_bits_iswrite),
    .io_MemResp_valid(WriteController_io_MemResp_valid),
    .io_MemResp_bits_data(WriteController_io_MemResp_bits_data),
    .io_MemResp_bits_tag(WriteController_io_MemResp_bits_tag)
  );
  ReadMemoryController ReadController ( // @[UnifiedController.scala 54:32]
    .clock(ReadController_clock),
    .reset(ReadController_reset),
    .io_ReadIn_0_ready(ReadController_io_ReadIn_0_ready),
    .io_ReadIn_0_valid(ReadController_io_ReadIn_0_valid),
    .io_ReadIn_0_bits_address(ReadController_io_ReadIn_0_bits_address),
    .io_ReadIn_0_bits_taskID(ReadController_io_ReadIn_0_bits_taskID),
    .io_ReadIn_1_ready(ReadController_io_ReadIn_1_ready),
    .io_ReadIn_1_valid(ReadController_io_ReadIn_1_valid),
    .io_ReadIn_1_bits_address(ReadController_io_ReadIn_1_bits_address),
    .io_ReadIn_1_bits_taskID(ReadController_io_ReadIn_1_bits_taskID),
    .io_ReadOut_0_valid(ReadController_io_ReadOut_0_valid),
    .io_ReadOut_0_data(ReadController_io_ReadOut_0_data),
    .io_ReadOut_1_valid(ReadController_io_ReadOut_1_valid),
    .io_ReadOut_1_data(ReadController_io_ReadOut_1_data),
    .io_MemReq_ready(ReadController_io_MemReq_ready),
    .io_MemReq_valid(ReadController_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadController_io_MemReq_bits_addr),
    .io_MemReq_bits_data(ReadController_io_MemReq_bits_data),
    .io_MemReq_bits_mask(ReadController_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(ReadController_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadController_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadController_io_MemReq_bits_iswrite),
    .io_MemResp_valid(ReadController_io_MemResp_valid),
    .io_MemResp_bits_data(ReadController_io_MemResp_bits_data),
    .io_MemResp_bits_tag(ReadController_io_MemResp_bits_tag)
  );
  ReadWriteArbiter ReadWriteArbiter ( // @[UnifiedController.scala 55:32]
    .clock(ReadWriteArbiter_clock),
    .io_ReadMemReq_ready(ReadWriteArbiter_io_ReadMemReq_ready),
    .io_ReadMemReq_valid(ReadWriteArbiter_io_ReadMemReq_valid),
    .io_ReadMemReq_bits_addr(ReadWriteArbiter_io_ReadMemReq_bits_addr),
    .io_ReadMemReq_bits_data(ReadWriteArbiter_io_ReadMemReq_bits_data),
    .io_ReadMemReq_bits_mask(ReadWriteArbiter_io_ReadMemReq_bits_mask),
    .io_ReadMemReq_bits_tag(ReadWriteArbiter_io_ReadMemReq_bits_tag),
    .io_ReadMemReq_bits_taskID(ReadWriteArbiter_io_ReadMemReq_bits_taskID),
    .io_ReadMemReq_bits_iswrite(ReadWriteArbiter_io_ReadMemReq_bits_iswrite),
    .io_WriteMemReq_ready(ReadWriteArbiter_io_WriteMemReq_ready),
    .io_WriteMemReq_valid(ReadWriteArbiter_io_WriteMemReq_valid),
    .io_WriteMemReq_bits_addr(ReadWriteArbiter_io_WriteMemReq_bits_addr),
    .io_WriteMemReq_bits_data(ReadWriteArbiter_io_WriteMemReq_bits_data),
    .io_WriteMemReq_bits_mask(ReadWriteArbiter_io_WriteMemReq_bits_mask),
    .io_WriteMemReq_bits_tag(ReadWriteArbiter_io_WriteMemReq_bits_tag),
    .io_WriteMemReq_bits_taskID(ReadWriteArbiter_io_WriteMemReq_bits_taskID),
    .io_WriteMemReq_bits_iswrite(ReadWriteArbiter_io_WriteMemReq_bits_iswrite),
    .io_MemResp_valid(ReadWriteArbiter_io_MemResp_valid),
    .io_MemResp_bits_data(ReadWriteArbiter_io_MemResp_bits_data),
    .io_MemResp_bits_tag(ReadWriteArbiter_io_MemResp_bits_tag),
    .io_MemResp_bits_iswrite(ReadWriteArbiter_io_MemResp_bits_iswrite),
    .io_ReadMemResp_valid(ReadWriteArbiter_io_ReadMemResp_valid),
    .io_ReadMemResp_bits_data(ReadWriteArbiter_io_ReadMemResp_bits_data),
    .io_ReadMemResp_bits_tag(ReadWriteArbiter_io_ReadMemResp_bits_tag),
    .io_WriteMemResp_valid(ReadWriteArbiter_io_WriteMemResp_valid),
    .io_WriteMemResp_bits_data(ReadWriteArbiter_io_WriteMemResp_bits_data),
    .io_WriteMemResp_bits_tag(ReadWriteArbiter_io_WriteMemResp_bits_tag),
    .io_MemReq_ready(ReadWriteArbiter_io_MemReq_ready),
    .io_MemReq_valid(ReadWriteArbiter_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadWriteArbiter_io_MemReq_bits_addr),
    .io_MemReq_bits_data(ReadWriteArbiter_io_MemReq_bits_data),
    .io_MemReq_bits_mask(ReadWriteArbiter_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(ReadWriteArbiter_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadWriteArbiter_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadWriteArbiter_io_MemReq_bits_iswrite)
  );
  assign _T = io_MemReq_ready & io_MemReq_valid; // @[Decoupled.scala 40:37]
  assign _T_1 = $unsigned(reset); // @[UnifiedController.scala 92:15]
  assign _T_2 = _T_1 == 1'h0; // @[UnifiedController.scala 92:15]
  assign io_WriteIn_0_ready = WriteController_io_WriteIn_0_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteOut_0_valid = WriteController_io_WriteOut_0_valid; // @[UnifiedController.scala 64:20]
  assign io_ReadIn_0_ready = ReadController_io_ReadIn_0_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_1_ready = ReadController_io_ReadIn_1_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadOut_0_valid = ReadController_io_ReadOut_0_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_0_data = ReadController_io_ReadOut_0_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_1_valid = ReadController_io_ReadOut_1_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_1_data = ReadController_io_ReadOut_1_data; // @[UnifiedController.scala 70:19]
  assign io_MemReq_valid = ReadWriteArbiter_io_MemReq_valid; // @[UnifiedController.scala 83:19]
  assign io_MemReq_bits_addr = ReadWriteArbiter_io_MemReq_bits_addr; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_data = ReadWriteArbiter_io_MemReq_bits_data; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_mask = ReadWriteArbiter_io_MemReq_bits_mask; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_tag = ReadWriteArbiter_io_MemReq_bits_tag; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_taskID = ReadWriteArbiter_io_MemReq_bits_taskID; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_iswrite = ReadWriteArbiter_io_MemReq_bits_iswrite; // @[UnifiedController.scala 82:18]
  assign WriteController_clock = clock;
  assign WriteController_reset = reset;
  assign WriteController_io_WriteIn_0_valid = io_WriteIn_0_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_0_bits_address = io_WriteIn_0_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_0_bits_data = io_WriteIn_0_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_0_bits_taskID = io_WriteIn_0_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_MemReq_ready = ReadWriteArbiter_io_WriteMemReq_ready; // @[UnifiedController.scala 77:35]
  assign WriteController_io_MemResp_valid = ReadWriteArbiter_io_WriteMemResp_valid; // @[UnifiedController.scala 78:30]
  assign WriteController_io_MemResp_bits_data = ReadWriteArbiter_io_WriteMemResp_bits_data; // @[UnifiedController.scala 78:30]
  assign WriteController_io_MemResp_bits_tag = ReadWriteArbiter_io_WriteMemResp_bits_tag; // @[UnifiedController.scala 78:30]
  assign ReadController_clock = clock;
  assign ReadController_reset = reset;
  assign ReadController_io_ReadIn_0_valid = io_ReadIn_0_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_0_bits_address = io_ReadIn_0_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_0_bits_taskID = io_ReadIn_0_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_1_valid = io_ReadIn_1_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_1_bits_address = io_ReadIn_1_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_1_bits_taskID = io_ReadIn_1_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_MemReq_ready = ReadWriteArbiter_io_ReadMemReq_ready; // @[UnifiedController.scala 74:34]
  assign ReadController_io_MemResp_valid = ReadWriteArbiter_io_ReadMemResp_valid; // @[UnifiedController.scala 75:29]
  assign ReadController_io_MemResp_bits_data = ReadWriteArbiter_io_ReadMemResp_bits_data; // @[UnifiedController.scala 75:29]
  assign ReadController_io_MemResp_bits_tag = ReadWriteArbiter_io_ReadMemResp_bits_tag; // @[UnifiedController.scala 75:29]
  assign ReadWriteArbiter_clock = clock;
  assign ReadWriteArbiter_io_ReadMemReq_valid = ReadController_io_MemReq_valid; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_addr = ReadController_io_MemReq_bits_addr; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_data = ReadController_io_MemReq_bits_data; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_mask = ReadController_io_MemReq_bits_mask; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_tag = ReadController_io_MemReq_bits_tag; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_taskID = ReadController_io_MemReq_bits_taskID; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_iswrite = ReadController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_WriteMemReq_valid = WriteController_io_MemReq_valid; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_addr = WriteController_io_MemReq_bits_addr; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_data = WriteController_io_MemReq_bits_data; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_mask = WriteController_io_MemReq_bits_mask; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_tag = WriteController_io_MemReq_bits_tag; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_taskID = WriteController_io_MemReq_bits_taskID; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_iswrite = WriteController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_MemResp_valid = io_MemResp_valid; // @[UnifiedController.scala 84:31]
  assign ReadWriteArbiter_io_MemResp_bits_data = io_MemResp_bits_data; // @[UnifiedController.scala 84:31]
  assign ReadWriteArbiter_io_MemResp_bits_tag = io_MemResp_bits_tag; // @[UnifiedController.scala 84:31]
  assign ReadWriteArbiter_io_MemResp_bits_iswrite = io_MemResp_bits_iswrite; // @[UnifiedController.scala 84:31]
  assign ReadWriteArbiter_io_MemReq_ready = io_MemReq_ready; // @[UnifiedController.scala 81:36]
  assign _GEN_0 = _T & io_MemReq_bits_iswrite; // @[UnifiedController.scala 92:15]
  assign _GEN_1 = io_MemReq_bits_iswrite == 1'h0; // @[UnifiedController.scala 94:15]
  assign _GEN_2 = _T & _GEN_1; // @[UnifiedController.scala 94:15]
  assign _GEN_3 = io_MemResp_valid & io_MemResp_bits_iswrite; // @[UnifiedController.scala 100:15]
  assign _GEN_4 = io_MemResp_bits_iswrite == 1'h0; // @[UnifiedController.scala 102:15]
  assign _GEN_5 = io_MemResp_valid & _GEN_4; // @[UnifiedController.scala 102:15]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_0 & _T_2) begin
          $fwrite(32'h80000002,"[LOG] [MemController] [MemReq]: Addr: %d, Data: %d, IsWrite: ST\n",io_MemReq_bits_addr,io_MemReq_bits_data); // @[UnifiedController.scala 92:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2 & _T_2) begin
          $fwrite(32'h80000002,"[LOG] [MemController] [MemReq]: Addr: %d, Data: %d, IsWrite: LD\n",io_MemReq_bits_addr,io_MemReq_bits_data); // @[UnifiedController.scala 94:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_3 & _T_2) begin
          $fwrite(32'h80000002,"[LOG] [MemController] [MemResp]: Data: %d, IsWrite: ST\n",io_MemResp_bits_data); // @[UnifiedController.scala 100:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & _T_2) begin
          $fwrite(32'h80000002,"[LOG] [MemController] [MemResp]: Data: %d, IsWrite: LD\n",io_MemReq_bits_data); // @[UnifiedController.scala 102:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SplitCallNew(
  input         clock,
  input         reset,
  output        io_In_ready,
  input         io_In_valid,
  input  [4:0]  io_In_bits_enable_taskID,
  input         io_In_bits_enable_control,
  input  [31:0] io_In_bits_data_field10_data,
  input  [31:0] io_In_bits_data_field9_data,
  input  [4:0]  io_In_bits_data_field8_taskID,
  input  [31:0] io_In_bits_data_field8_data,
  input  [31:0] io_In_bits_data_field7_data,
  input  [4:0]  io_In_bits_data_field6_taskID,
  input  [31:0] io_In_bits_data_field6_data,
  input  [31:0] io_In_bits_data_field5_data,
  input  [4:0]  io_In_bits_data_field4_taskID,
  input  [31:0] io_In_bits_data_field4_data,
  input  [31:0] io_In_bits_data_field3_data,
  input  [31:0] io_In_bits_data_field2_data,
  input  [4:0]  io_In_bits_data_field1_taskID,
  input  [31:0] io_In_bits_data_field1_data,
  input  [4:0]  io_In_bits_data_field0_taskID,
  input  [31:0] io_In_bits_data_field0_data,
  input         io_Out_enable_ready,
  output        io_Out_enable_valid,
  output [4:0]  io_Out_enable_bits_taskID,
  output        io_Out_enable_bits_control,
  input         io_Out_data_field10_0_ready,
  output        io_Out_data_field10_0_valid,
  output [31:0] io_Out_data_field10_0_bits_data,
  input         io_Out_data_field9_0_ready,
  output        io_Out_data_field9_0_valid,
  output [31:0] io_Out_data_field9_0_bits_data,
  input         io_Out_data_field8_0_ready,
  output        io_Out_data_field8_0_valid,
  output [4:0]  io_Out_data_field8_0_bits_taskID,
  output [31:0] io_Out_data_field8_0_bits_data,
  input         io_Out_data_field8_1_ready,
  output        io_Out_data_field8_1_valid,
  output [31:0] io_Out_data_field8_1_bits_data,
  input         io_Out_data_field8_2_ready,
  output        io_Out_data_field8_2_valid,
  output [31:0] io_Out_data_field8_2_bits_data,
  input         io_Out_data_field7_0_ready,
  output        io_Out_data_field7_0_valid,
  output [31:0] io_Out_data_field7_0_bits_data,
  input         io_Out_data_field7_1_ready,
  output        io_Out_data_field7_1_valid,
  output [31:0] io_Out_data_field7_1_bits_data,
  input         io_Out_data_field6_0_ready,
  output        io_Out_data_field6_0_valid,
  output [4:0]  io_Out_data_field6_0_bits_taskID,
  output [31:0] io_Out_data_field6_0_bits_data,
  input         io_Out_data_field6_1_ready,
  output        io_Out_data_field6_1_valid,
  output [31:0] io_Out_data_field6_1_bits_data,
  input         io_Out_data_field6_2_ready,
  output        io_Out_data_field6_2_valid,
  output [31:0] io_Out_data_field6_2_bits_data,
  input         io_Out_data_field5_0_ready,
  output        io_Out_data_field5_0_valid,
  output [31:0] io_Out_data_field5_0_bits_data,
  input         io_Out_data_field5_1_ready,
  output        io_Out_data_field5_1_valid,
  output [31:0] io_Out_data_field5_1_bits_data,
  input         io_Out_data_field4_0_ready,
  output        io_Out_data_field4_0_valid,
  output [4:0]  io_Out_data_field4_0_bits_taskID,
  output [31:0] io_Out_data_field4_0_bits_data,
  input         io_Out_data_field4_1_ready,
  output        io_Out_data_field4_1_valid,
  output [31:0] io_Out_data_field4_1_bits_data,
  input         io_Out_data_field4_2_ready,
  output        io_Out_data_field4_2_valid,
  output [31:0] io_Out_data_field4_2_bits_data,
  input         io_Out_data_field3_0_ready,
  output        io_Out_data_field3_0_valid,
  output [31:0] io_Out_data_field3_0_bits_data,
  input         io_Out_data_field2_0_ready,
  output        io_Out_data_field2_0_valid,
  output [31:0] io_Out_data_field2_0_bits_data,
  input         io_Out_data_field1_0_ready,
  output        io_Out_data_field1_0_valid,
  output [4:0]  io_Out_data_field1_0_bits_taskID,
  output [31:0] io_Out_data_field1_0_bits_data,
  input         io_Out_data_field0_0_ready,
  output        io_Out_data_field0_0_valid,
  output [4:0]  io_Out_data_field0_0_bits_taskID,
  output [31:0] io_Out_data_field0_0_bits_data
);
  reg [4:0] inputReg_enable_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_0;
  reg  inputReg_enable_control; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_1;
  reg [31:0] inputReg_data_field10_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_2;
  reg [31:0] inputReg_data_field9_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_3;
  reg [4:0] inputReg_data_field8_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_4;
  reg [31:0] inputReg_data_field8_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_5;
  reg [31:0] inputReg_data_field7_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_6;
  reg [4:0] inputReg_data_field6_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_7;
  reg [31:0] inputReg_data_field6_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_8;
  reg [31:0] inputReg_data_field5_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_9;
  reg [4:0] inputReg_data_field4_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_10;
  reg [31:0] inputReg_data_field4_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_11;
  reg [31:0] inputReg_data_field3_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_12;
  reg [31:0] inputReg_data_field2_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_13;
  reg [4:0] inputReg_data_field1_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_14;
  reg [31:0] inputReg_data_field1_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_15;
  reg [4:0] inputReg_data_field0_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_16;
  reg [31:0] inputReg_data_field0_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_17;
  reg  enableValidReg; // @[SplitDecoupled.scala 154:31]
  reg [31:0] _RAND_18;
  reg  allValid_0; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_19;
  reg  allValid_1; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_20;
  reg  allValid_2; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_21;
  reg  allValid_3; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_22;
  reg  outputValidReg_4_0; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_23;
  reg  outputValidReg_4_1; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_24;
  reg  outputValidReg_4_2; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_25;
  reg  outputValidReg_5_0; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_26;
  reg  outputValidReg_5_1; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_27;
  reg  outputValidReg_6_0; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_28;
  reg  outputValidReg_6_1; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_29;
  reg  outputValidReg_6_2; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_30;
  reg  outputValidReg_7_0; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_31;
  reg  outputValidReg_7_1; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_32;
  reg  outputValidReg_8_0; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_33;
  reg  outputValidReg_8_1; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_34;
  reg  outputValidReg_8_2; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_35;
  reg  allValid_9; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_36;
  reg  allValid_10; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_37;
  wire  _T_37; // @[SplitDecoupled.scala 161:51]
  wire  allValid_4; // @[SplitDecoupled.scala 161:51]
  wire  allValid_5; // @[SplitDecoupled.scala 161:51]
  wire  _T_38; // @[SplitDecoupled.scala 161:51]
  wire  allValid_6; // @[SplitDecoupled.scala 161:51]
  wire  allValid_7; // @[SplitDecoupled.scala 161:51]
  wire  _T_39; // @[SplitDecoupled.scala 161:51]
  wire  allValid_8; // @[SplitDecoupled.scala 161:51]
  reg  state; // @[SplitDecoupled.scala 166:22]
  reg [31:0] _RAND_38;
  wire  _T_40; // @[SplitDecoupled.scala 168:24]
  wire  _T_41; // @[Conditional.scala 37:30]
  wire  _T_42; // @[Decoupled.scala 40:37]
  wire  _GEN_0; // @[SplitDecoupled.scala 172:27]
  wire  _T_44; // @[SplitDecoupled.scala 178:36]
  wire  _T_45; // @[SplitDecoupled.scala 178:36]
  wire  _T_46; // @[SplitDecoupled.scala 178:36]
  wire  _T_47; // @[SplitDecoupled.scala 178:36]
  wire  _T_48; // @[SplitDecoupled.scala 178:36]
  wire  _T_49; // @[SplitDecoupled.scala 178:36]
  wire  _T_50; // @[SplitDecoupled.scala 178:36]
  wire  _T_51; // @[SplitDecoupled.scala 178:36]
  wire  _T_52; // @[SplitDecoupled.scala 178:36]
  wire  _T_53; // @[SplitDecoupled.scala 178:36]
  wire  _T_54; // @[SplitDecoupled.scala 178:13]
  wire  _T_55; // @[SplitDecoupled.scala 178:45]
  wire  _T_56; // @[SplitDecoupled.scala 178:42]
  wire  _T_58; // @[SplitDecoupled.scala 186:24]
  wire  _GEN_74; // @[SplitDecoupled.scala 186:45]
  wire  _T_60; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_76; // @[SplitDecoupled.scala 186:45]
  wire  _T_64; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_78; // @[SplitDecoupled.scala 186:45]
  wire  _T_68; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_80; // @[SplitDecoupled.scala 186:45]
  wire  _T_72; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_82; // @[SplitDecoupled.scala 186:45]
  wire  _T_76; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_84; // @[SplitDecoupled.scala 186:45]
  wire  _T_80; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_86; // @[SplitDecoupled.scala 186:45]
  wire  _T_84; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_88; // @[SplitDecoupled.scala 186:45]
  wire  _T_88; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_90; // @[SplitDecoupled.scala 186:45]
  wire  _T_92; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_92; // @[SplitDecoupled.scala 186:45]
  wire  _T_96; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_94; // @[SplitDecoupled.scala 186:45]
  wire  _T_100; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_96; // @[SplitDecoupled.scala 186:45]
  wire  _T_104; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_98; // @[SplitDecoupled.scala 186:45]
  wire  _T_108; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_100; // @[SplitDecoupled.scala 186:45]
  wire  _T_112; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_102; // @[SplitDecoupled.scala 186:45]
  wire  _T_116; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_104; // @[SplitDecoupled.scala 186:45]
  wire  _T_120; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_106; // @[SplitDecoupled.scala 186:45]
  wire  _T_124; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_108; // @[SplitDecoupled.scala 186:45]
  wire  _T_128; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_110; // @[SplitDecoupled.scala 186:45]
  wire  _T_132; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_112; // @[SplitDecoupled.scala 197:41]
  wire  _T_136; // @[SplitDecoupled.scala 200:28]
  assign _T_37 = outputValidReg_4_0 | outputValidReg_4_1; // @[SplitDecoupled.scala 161:51]
  assign allValid_4 = _T_37 | outputValidReg_4_2; // @[SplitDecoupled.scala 161:51]
  assign allValid_5 = outputValidReg_5_0 | outputValidReg_5_1; // @[SplitDecoupled.scala 161:51]
  assign _T_38 = outputValidReg_6_0 | outputValidReg_6_1; // @[SplitDecoupled.scala 161:51]
  assign allValid_6 = _T_38 | outputValidReg_6_2; // @[SplitDecoupled.scala 161:51]
  assign allValid_7 = outputValidReg_7_0 | outputValidReg_7_1; // @[SplitDecoupled.scala 161:51]
  assign _T_39 = outputValidReg_8_0 | outputValidReg_8_1; // @[SplitDecoupled.scala 161:51]
  assign allValid_8 = _T_39 | outputValidReg_8_2; // @[SplitDecoupled.scala 161:51]
  assign _T_40 = state == 1'h0; // @[SplitDecoupled.scala 168:24]
  assign _T_41 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_42 = io_In_ready & io_In_valid; // @[Decoupled.scala 40:37]
  assign _GEN_0 = _T_42 | state; // @[SplitDecoupled.scala 172:27]
  assign _T_44 = allValid_0 | allValid_1; // @[SplitDecoupled.scala 178:36]
  assign _T_45 = _T_44 | allValid_2; // @[SplitDecoupled.scala 178:36]
  assign _T_46 = _T_45 | allValid_3; // @[SplitDecoupled.scala 178:36]
  assign _T_47 = _T_46 | allValid_4; // @[SplitDecoupled.scala 178:36]
  assign _T_48 = _T_47 | allValid_5; // @[SplitDecoupled.scala 178:36]
  assign _T_49 = _T_48 | allValid_6; // @[SplitDecoupled.scala 178:36]
  assign _T_50 = _T_49 | allValid_7; // @[SplitDecoupled.scala 178:36]
  assign _T_51 = _T_50 | allValid_8; // @[SplitDecoupled.scala 178:36]
  assign _T_52 = _T_51 | allValid_9; // @[SplitDecoupled.scala 178:36]
  assign _T_53 = _T_52 | allValid_10; // @[SplitDecoupled.scala 178:36]
  assign _T_54 = _T_53 == 1'h0; // @[SplitDecoupled.scala 178:13]
  assign _T_55 = enableValidReg == 1'h0; // @[SplitDecoupled.scala 178:45]
  assign _T_56 = _T_54 & _T_55; // @[SplitDecoupled.scala 178:42]
  assign _T_58 = io_In_valid & _T_40; // @[SplitDecoupled.scala 186:24]
  assign _GEN_74 = _T_58 | allValid_0; // @[SplitDecoupled.scala 186:45]
  assign _T_60 = state & io_Out_data_field0_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_76 = _T_58 | allValid_1; // @[SplitDecoupled.scala 186:45]
  assign _T_64 = state & io_Out_data_field1_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_78 = _T_58 | allValid_2; // @[SplitDecoupled.scala 186:45]
  assign _T_68 = state & io_Out_data_field2_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_80 = _T_58 | allValid_3; // @[SplitDecoupled.scala 186:45]
  assign _T_72 = state & io_Out_data_field3_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_82 = _T_58 | outputValidReg_4_0; // @[SplitDecoupled.scala 186:45]
  assign _T_76 = state & io_Out_data_field4_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_84 = _T_58 | outputValidReg_4_1; // @[SplitDecoupled.scala 186:45]
  assign _T_80 = state & io_Out_data_field4_1_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_86 = _T_58 | outputValidReg_4_2; // @[SplitDecoupled.scala 186:45]
  assign _T_84 = state & io_Out_data_field4_2_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_88 = _T_58 | outputValidReg_5_0; // @[SplitDecoupled.scala 186:45]
  assign _T_88 = state & io_Out_data_field5_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_90 = _T_58 | outputValidReg_5_1; // @[SplitDecoupled.scala 186:45]
  assign _T_92 = state & io_Out_data_field5_1_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_92 = _T_58 | outputValidReg_6_0; // @[SplitDecoupled.scala 186:45]
  assign _T_96 = state & io_Out_data_field6_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_94 = _T_58 | outputValidReg_6_1; // @[SplitDecoupled.scala 186:45]
  assign _T_100 = state & io_Out_data_field6_1_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_96 = _T_58 | outputValidReg_6_2; // @[SplitDecoupled.scala 186:45]
  assign _T_104 = state & io_Out_data_field6_2_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_98 = _T_58 | outputValidReg_7_0; // @[SplitDecoupled.scala 186:45]
  assign _T_108 = state & io_Out_data_field7_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_100 = _T_58 | outputValidReg_7_1; // @[SplitDecoupled.scala 186:45]
  assign _T_112 = state & io_Out_data_field7_1_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_102 = _T_58 | outputValidReg_8_0; // @[SplitDecoupled.scala 186:45]
  assign _T_116 = state & io_Out_data_field8_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_104 = _T_58 | outputValidReg_8_1; // @[SplitDecoupled.scala 186:45]
  assign _T_120 = state & io_Out_data_field8_1_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_106 = _T_58 | outputValidReg_8_2; // @[SplitDecoupled.scala 186:45]
  assign _T_124 = state & io_Out_data_field8_2_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_108 = _T_58 | allValid_9; // @[SplitDecoupled.scala 186:45]
  assign _T_128 = state & io_Out_data_field9_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_110 = _T_58 | allValid_10; // @[SplitDecoupled.scala 186:45]
  assign _T_132 = state & io_Out_data_field10_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_112 = _T_58 | enableValidReg; // @[SplitDecoupled.scala 197:41]
  assign _T_136 = state & io_Out_enable_ready; // @[SplitDecoupled.scala 200:28]
  assign io_In_ready = state == 1'h0; // @[SplitDecoupled.scala 168:15]
  assign io_Out_enable_valid = enableValidReg; // @[SplitDecoupled.scala 203:23]
  assign io_Out_enable_bits_taskID = inputReg_enable_taskID; // @[SplitDecoupled.scala 204:22]
  assign io_Out_enable_bits_control = inputReg_enable_control; // @[SplitDecoupled.scala 204:22]
  assign io_Out_data_field10_0_valid = allValid_10; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field10_0_bits_data = inputReg_data_field10_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field9_0_valid = allValid_9; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field9_0_bits_data = inputReg_data_field9_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field8_0_valid = outputValidReg_8_0; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field8_0_bits_taskID = inputReg_data_field8_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field8_0_bits_data = inputReg_data_field8_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field8_1_valid = outputValidReg_8_1; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field8_1_bits_data = inputReg_data_field8_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field8_2_valid = outputValidReg_8_2; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field8_2_bits_data = inputReg_data_field8_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field7_0_valid = outputValidReg_7_0; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field7_0_bits_data = inputReg_data_field7_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field7_1_valid = outputValidReg_7_1; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field7_1_bits_data = inputReg_data_field7_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field6_0_valid = outputValidReg_6_0; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field6_0_bits_taskID = inputReg_data_field6_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field6_0_bits_data = inputReg_data_field6_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field6_1_valid = outputValidReg_6_1; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field6_1_bits_data = inputReg_data_field6_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field6_2_valid = outputValidReg_6_2; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field6_2_bits_data = inputReg_data_field6_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field5_0_valid = outputValidReg_5_0; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field5_0_bits_data = inputReg_data_field5_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field5_1_valid = outputValidReg_5_1; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field5_1_bits_data = inputReg_data_field5_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field4_0_valid = outputValidReg_4_0; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field4_0_bits_taskID = inputReg_data_field4_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field4_0_bits_data = inputReg_data_field4_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field4_1_valid = outputValidReg_4_1; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field4_1_bits_data = inputReg_data_field4_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field4_2_valid = outputValidReg_4_2; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field4_2_bits_data = inputReg_data_field4_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field3_0_valid = allValid_3; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field3_0_bits_data = inputReg_data_field3_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field2_0_valid = allValid_2; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field2_0_bits_data = inputReg_data_field2_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_0_valid = allValid_1; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_0_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_0_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field0_0_valid = allValid_0; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field0_0_bits_taskID = inputReg_data_field0_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field0_0_bits_data = inputReg_data_field0_data; // @[SplitDecoupled.scala 193:39]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inputReg_enable_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inputReg_enable_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inputReg_data_field10_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  inputReg_data_field9_data = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  inputReg_data_field8_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  inputReg_data_field8_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  inputReg_data_field7_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inputReg_data_field6_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  inputReg_data_field6_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  inputReg_data_field5_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  inputReg_data_field4_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  inputReg_data_field4_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  inputReg_data_field3_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  inputReg_data_field2_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  inputReg_data_field1_taskID = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  inputReg_data_field1_data = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  inputReg_data_field0_taskID = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  inputReg_data_field0_data = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  enableValidReg = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  allValid_0 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  allValid_1 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  allValid_2 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  allValid_3 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  outputValidReg_4_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  outputValidReg_4_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  outputValidReg_4_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  outputValidReg_5_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  outputValidReg_5_1 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  outputValidReg_6_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  outputValidReg_6_1 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  outputValidReg_6_2 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  outputValidReg_7_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  outputValidReg_7_1 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  outputValidReg_8_0 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  outputValidReg_8_1 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  outputValidReg_8_2 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  allValid_9 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  allValid_10 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  state = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      inputReg_enable_taskID <= 5'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_enable_taskID <= io_In_bits_enable_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_enable_control <= 1'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_enable_control <= io_In_bits_enable_control;
        end
      end
    end
    if (reset) begin
      inputReg_data_field10_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field10_data <= io_In_bits_data_field10_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field9_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field9_data <= io_In_bits_data_field9_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field8_taskID <= 5'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field8_taskID <= io_In_bits_data_field8_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field8_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field8_data <= io_In_bits_data_field8_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field7_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field7_data <= io_In_bits_data_field7_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field6_taskID <= 5'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field6_taskID <= io_In_bits_data_field6_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field6_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field6_data <= io_In_bits_data_field6_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field5_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field5_data <= io_In_bits_data_field5_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field4_taskID <= 5'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field4_taskID <= io_In_bits_data_field4_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field4_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field4_data <= io_In_bits_data_field4_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field3_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field3_data <= io_In_bits_data_field3_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field2_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field2_data <= io_In_bits_data_field2_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field1_taskID <= 5'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field1_taskID <= io_In_bits_data_field1_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field1_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field1_data <= io_In_bits_data_field1_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field0_taskID <= 5'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field0_taskID <= io_In_bits_data_field0_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field0_data <= 32'h0;
    end else begin
      if (_T_41) begin
        if (_T_42) begin
          inputReg_data_field0_data <= io_In_bits_data_field0_data;
        end
      end
    end
    if (reset) begin
      enableValidReg <= 1'h0;
    end else begin
      if (_T_136) begin
        enableValidReg <= 1'h0;
      end else begin
        enableValidReg <= _GEN_112;
      end
    end
    if (reset) begin
      allValid_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        allValid_0 <= 1'h0;
      end else begin
        allValid_0 <= _GEN_74;
      end
    end
    if (reset) begin
      allValid_1 <= 1'h0;
    end else begin
      if (_T_64) begin
        allValid_1 <= 1'h0;
      end else begin
        allValid_1 <= _GEN_76;
      end
    end
    if (reset) begin
      allValid_2 <= 1'h0;
    end else begin
      if (_T_68) begin
        allValid_2 <= 1'h0;
      end else begin
        allValid_2 <= _GEN_78;
      end
    end
    if (reset) begin
      allValid_3 <= 1'h0;
    end else begin
      if (_T_72) begin
        allValid_3 <= 1'h0;
      end else begin
        allValid_3 <= _GEN_80;
      end
    end
    if (reset) begin
      outputValidReg_4_0 <= 1'h0;
    end else begin
      if (_T_76) begin
        outputValidReg_4_0 <= 1'h0;
      end else begin
        outputValidReg_4_0 <= _GEN_82;
      end
    end
    if (reset) begin
      outputValidReg_4_1 <= 1'h0;
    end else begin
      if (_T_80) begin
        outputValidReg_4_1 <= 1'h0;
      end else begin
        outputValidReg_4_1 <= _GEN_84;
      end
    end
    if (reset) begin
      outputValidReg_4_2 <= 1'h0;
    end else begin
      if (_T_84) begin
        outputValidReg_4_2 <= 1'h0;
      end else begin
        outputValidReg_4_2 <= _GEN_86;
      end
    end
    if (reset) begin
      outputValidReg_5_0 <= 1'h0;
    end else begin
      if (_T_88) begin
        outputValidReg_5_0 <= 1'h0;
      end else begin
        outputValidReg_5_0 <= _GEN_88;
      end
    end
    if (reset) begin
      outputValidReg_5_1 <= 1'h0;
    end else begin
      if (_T_92) begin
        outputValidReg_5_1 <= 1'h0;
      end else begin
        outputValidReg_5_1 <= _GEN_90;
      end
    end
    if (reset) begin
      outputValidReg_6_0 <= 1'h0;
    end else begin
      if (_T_96) begin
        outputValidReg_6_0 <= 1'h0;
      end else begin
        outputValidReg_6_0 <= _GEN_92;
      end
    end
    if (reset) begin
      outputValidReg_6_1 <= 1'h0;
    end else begin
      if (_T_100) begin
        outputValidReg_6_1 <= 1'h0;
      end else begin
        outputValidReg_6_1 <= _GEN_94;
      end
    end
    if (reset) begin
      outputValidReg_6_2 <= 1'h0;
    end else begin
      if (_T_104) begin
        outputValidReg_6_2 <= 1'h0;
      end else begin
        outputValidReg_6_2 <= _GEN_96;
      end
    end
    if (reset) begin
      outputValidReg_7_0 <= 1'h0;
    end else begin
      if (_T_108) begin
        outputValidReg_7_0 <= 1'h0;
      end else begin
        outputValidReg_7_0 <= _GEN_98;
      end
    end
    if (reset) begin
      outputValidReg_7_1 <= 1'h0;
    end else begin
      if (_T_112) begin
        outputValidReg_7_1 <= 1'h0;
      end else begin
        outputValidReg_7_1 <= _GEN_100;
      end
    end
    if (reset) begin
      outputValidReg_8_0 <= 1'h0;
    end else begin
      if (_T_116) begin
        outputValidReg_8_0 <= 1'h0;
      end else begin
        outputValidReg_8_0 <= _GEN_102;
      end
    end
    if (reset) begin
      outputValidReg_8_1 <= 1'h0;
    end else begin
      if (_T_120) begin
        outputValidReg_8_1 <= 1'h0;
      end else begin
        outputValidReg_8_1 <= _GEN_104;
      end
    end
    if (reset) begin
      outputValidReg_8_2 <= 1'h0;
    end else begin
      if (_T_124) begin
        outputValidReg_8_2 <= 1'h0;
      end else begin
        outputValidReg_8_2 <= _GEN_106;
      end
    end
    if (reset) begin
      allValid_9 <= 1'h0;
    end else begin
      if (_T_128) begin
        allValid_9 <= 1'h0;
      end else begin
        allValid_9 <= _GEN_108;
      end
    end
    if (reset) begin
      allValid_10 <= 1'h0;
    end else begin
      if (_T_132) begin
        allValid_10 <= 1'h0;
      end else begin
        allValid_10 <= _GEN_110;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_41) begin
        state <= _GEN_0;
      end else begin
        if (state) begin
          if (_T_56) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module LoopBlockNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [4:0]  io_InLiveIn_0_bits_taskID,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [4:0]  io_InLiveIn_2_bits_taskID,
  input  [31:0] io_InLiveIn_2_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [4:0]  io_OutLiveIn_field2_0_bits_taskID,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [4:0]  io_OutLiveIn_field0_0_bits_taskID,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  output        io_CarryDepenIn_1_ready,
  input         io_CarryDepenIn_1_valid,
  input  [4:0]  io_CarryDepenIn_1_bits_taskID,
  input  [31:0] io_CarryDepenIn_1_bits_data,
  input         io_CarryDepenOut_field1_0_ready,
  output        io_CarryDepenOut_field1_0_valid,
  output [4:0]  io_CarryDepenOut_field1_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field1_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  output        io_InLiveOut_0_ready,
  input         io_InLiveOut_0_valid,
  input  [4:0]  io_InLiveOut_0_bits_taskID,
  input  [31:0] io_InLiveOut_0_bits_data,
  input         io_OutLiveOut_field0_0_ready,
  output        io_OutLiveOut_field0_0_valid,
  output [4:0]  io_OutLiveOut_field0_0_bits_taskID,
  output [31:0] io_OutLiveOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_2;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_3;
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_5;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_6;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_7;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_8;
  reg [4:0] in_live_in_R_0_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [4:0] in_live_in_R_2_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_14;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_15;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_16;
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_17;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_18;
  reg [4:0] in_carry_in_R_1_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_19;
  reg [31:0] in_carry_in_R_1_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_20;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_21;
  reg  in_carry_in_valid_R_1; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_22;
  reg [4:0] in_live_out_R_0_taskID; // @[LoopBlock.scala 543:55]
  reg [31:0] _RAND_23;
  reg [31:0] in_live_out_R_0_data; // @[LoopBlock.scala 543:55]
  reg [31:0] _RAND_24;
  reg  in_live_out_valid_R_0; // @[LoopBlock.scala 544:61]
  reg [31:0] _RAND_25;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_26;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_27;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_28;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_29;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_30;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_31;
  reg  out_live_out_valid_R_0_0; // @[LoopBlock.scala 563:47]
  reg [31:0] _RAND_32;
  reg  out_live_out_fire_R_0_0; // @[LoopBlock.scala 567:47]
  reg [31:0] _RAND_33;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_34;
  reg  out_carry_out_valid_R_1_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_35;
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_36;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_37;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_38;
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_39;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_40;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_41;
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_42;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_43;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_44;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_45;
  wire  _T_17; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_19; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[LoopBlock.scala 603:33]
  wire [4:0] _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_25; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_27; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_29; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[LoopBlock.scala 632:34]
  wire  _T_31; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[LoopBlock.scala 641:37]
  wire  _T_33; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[LoopBlock.scala 641:37]
  wire  _T_34; // @[Decoupled.scala 40:37]
  wire  _GEN_34; // @[LoopBlock.scala 704:39]
  wire  _T_35; // @[Decoupled.scala 40:37]
  wire  _GEN_35; // @[LoopBlock.scala 708:38]
  wire  _T_36; // @[Decoupled.scala 40:37]
  wire  _GEN_36; // @[LoopBlock.scala 713:33]
  wire  _GEN_37; // @[LoopBlock.scala 713:33]
  wire  _T_37; // @[Decoupled.scala 40:37]
  wire  _GEN_38; // @[LoopBlock.scala 722:57]
  wire  _GEN_39; // @[LoopBlock.scala 722:57]
  wire  _T_38; // @[Decoupled.scala 40:37]
  wire  _GEN_40; // @[LoopBlock.scala 722:57]
  wire  _GEN_41; // @[LoopBlock.scala 722:57]
  wire  _T_39; // @[Decoupled.scala 40:37]
  wire  _GEN_42; // @[LoopBlock.scala 722:57]
  wire  _GEN_43; // @[LoopBlock.scala 722:57]
  wire  _T_40; // @[Decoupled.scala 40:37]
  wire  _GEN_44; // @[LoopBlock.scala 732:58]
  wire  _GEN_45; // @[LoopBlock.scala 732:58]
  wire  _T_41; // @[Decoupled.scala 40:37]
  wire  _GEN_46; // @[LoopBlock.scala 742:61]
  wire  _T_42; // @[Decoupled.scala 40:37]
  wire  _GEN_48; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_46;
  wire  _T_43; // @[Conditional.scala 37:30]
  wire  _T_44; // @[LoopBlock.scala 765:35]
  wire  _T_45; // @[LoopBlock.scala 765:35]
  wire  _T_46; // @[LoopBlock.scala 869:28]
  wire  _GEN_50; // @[LoopBlock.scala 870:26]
  wire  _GEN_51; // @[LoopBlock.scala 870:26]
  wire  _GEN_52; // @[LoopBlock.scala 870:26]
  wire  _GEN_53; // @[LoopBlock.scala 870:26]
  wire  _GEN_54; // @[LoopBlock.scala 870:26]
  wire  _GEN_55; // @[LoopBlock.scala 870:26]
  wire  _GEN_57; // @[LoopBlock.scala 870:26]
  wire  _GEN_60; // @[LoopBlock.scala 870:26]
  wire  _GEN_66; // @[LoopBlock.scala 870:26]
  wire  _T_51; // @[Conditional.scala 37:30]
  wire  _T_52; // @[LoopBlock.scala 898:30]
  wire  _T_53; // @[LoopBlock.scala 899:9]
  wire  _T_54; // @[LoopBlock.scala 828:26]
  wire  _T_55; // @[LoopBlock.scala 828:26]
  wire  _T_56; // @[LoopBlock.scala 899:29]
  wire  _T_57; // @[LoopBlock.scala 783:40]
  wire  _T_58; // @[LoopBlock.scala 900:9]
  wire  _T_64; // @[LoopBlock.scala 932:19]
  wire  _T_65; // @[LoopBlock.scala 932:19]
  wire  _GEN_88; // @[LoopBlock.scala 936:64]
  wire  _GEN_89; // @[LoopBlock.scala 936:64]
  wire  _GEN_92; // @[LoopBlock.scala 936:64]
  wire  _GEN_94; // @[LoopBlock.scala 936:64]
  wire  _GEN_99; // @[LoopBlock.scala 903:56]
  wire  _GEN_100; // @[LoopBlock.scala 903:56]
  wire  _GEN_102; // @[LoopBlock.scala 903:56]
  wire  _GEN_108; // @[LoopBlock.scala 903:56]
  wire  _GEN_109; // @[LoopBlock.scala 903:56]
  wire  _GEN_110; // @[LoopBlock.scala 903:56]
  wire  _GEN_111; // @[LoopBlock.scala 903:56]
  wire  _GEN_112; // @[LoopBlock.scala 903:56]
  wire  _T_75; // @[Conditional.scala 37:30]
  wire  _T_76; // @[LoopBlock.scala 963:27]
  wire  _GEN_300; // @[LoopBlock.scala 932:19]
  wire  _GEN_301; // @[LoopBlock.scala 932:19]
  wire  _GEN_302; // @[LoopBlock.scala 932:19]
  wire  _GEN_303; // @[LoopBlock.scala 932:19]
  wire  _GEN_307; // @[LoopBlock.scala 950:19]
  wire  _GEN_308; // @[LoopBlock.scala 950:19]
  wire  _GEN_309; // @[LoopBlock.scala 950:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_17 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_17 | enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_19 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_19 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_19 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_19 | loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_21 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_21 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_21 | loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_23 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_23 | in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_25 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_25 | in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_27 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_27 | in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_29 = io_InLiveOut_0_ready & io_InLiveOut_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_29 | in_live_out_valid_R_0; // @[LoopBlock.scala 632:34]
  assign _T_31 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_31 | in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_33 = io_CarryDepenIn_1_ready & io_CarryDepenIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_33 | in_carry_in_valid_R_1; // @[LoopBlock.scala 641:37]
  assign _T_34 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  assign _GEN_34 = _T_34 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_35 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  assign _GEN_35 = _T_35 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_36 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_36 = _T_36 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_37 = _T_36 | loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_37 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_38 = _T_37 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_39 = _T_37 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_38 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_40 = _T_38 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_41 = _T_38 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_39 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_42 = _T_39 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_43 = _T_39 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_40 = io_OutLiveOut_field0_0_ready & io_OutLiveOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_44 = _T_40 ? 1'h0 : out_live_out_valid_R_0_0; // @[LoopBlock.scala 732:58]
  assign _GEN_45 = _T_40 | out_live_out_fire_R_0_0; // @[LoopBlock.scala 732:58]
  assign _T_41 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_46 = _T_41 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_42 = io_CarryDepenOut_field1_0_ready & io_CarryDepenOut_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_48 = _T_42 ? 1'h0 : out_carry_out_valid_R_1_0; // @[LoopBlock.scala 742:61]
  assign _T_43 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_44 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_45 = _T_44 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_46 = _T_45 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_50 = enable_R_control | _GEN_38; // @[LoopBlock.scala 870:26]
  assign _GEN_51 = enable_R_control | _GEN_40; // @[LoopBlock.scala 870:26]
  assign _GEN_52 = enable_R_control | _GEN_42; // @[LoopBlock.scala 870:26]
  assign _GEN_53 = enable_R_control | _GEN_46; // @[LoopBlock.scala 870:26]
  assign _GEN_54 = enable_R_control | _GEN_48; // @[LoopBlock.scala 870:26]
  assign _GEN_55 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_57 = enable_R_control | _GEN_34; // @[LoopBlock.scala 870:26]
  assign _GEN_60 = enable_R_control | _GEN_35; // @[LoopBlock.scala 870:26]
  assign _GEN_66 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 870:26]
  assign _T_51 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_52 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_53 = _T_52 & in_live_out_valid_R_0; // @[LoopBlock.scala 899:9]
  assign _T_54 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_55 = _T_54 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_56 = _T_53 & _T_55; // @[LoopBlock.scala 899:29]
  assign _T_57 = in_carry_in_valid_R_0 & in_carry_in_valid_R_1; // @[LoopBlock.scala 783:40]
  assign _T_58 = _T_56 & _T_57; // @[LoopBlock.scala 900:9]
  assign _T_64 = $unsigned(reset); // @[LoopBlock.scala 932:19]
  assign _T_65 = _T_64 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_88 = loop_finish_R_0_control | _GEN_44; // @[LoopBlock.scala 936:64]
  assign _GEN_89 = loop_finish_R_0_control | _GEN_36; // @[LoopBlock.scala 936:64]
  assign _GEN_92 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_94 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_99 = loop_back_R_0_control | _GEN_34; // @[LoopBlock.scala 903:56]
  assign _GEN_100 = loop_back_R_0_control | _GEN_92; // @[LoopBlock.scala 903:56]
  assign _GEN_102 = loop_back_R_0_control | _GEN_35; // @[LoopBlock.scala 903:56]
  assign _GEN_108 = loop_back_R_0_control | _GEN_38; // @[LoopBlock.scala 903:56]
  assign _GEN_109 = loop_back_R_0_control | _GEN_40; // @[LoopBlock.scala 903:56]
  assign _GEN_110 = loop_back_R_0_control | _GEN_42; // @[LoopBlock.scala 903:56]
  assign _GEN_111 = loop_back_R_0_control | _GEN_46; // @[LoopBlock.scala 903:56]
  assign _GEN_112 = loop_back_R_0_control | _GEN_48; // @[LoopBlock.scala 903:56]
  assign _T_75 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_76 = loop_exit_fire_R_0 & out_live_out_fire_R_0_0; // @[LoopBlock.scala 963:27]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_taskID = in_live_in_R_2_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_taskID = in_live_in_R_0_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenIn_1_ready = ~ in_carry_in_valid_R_1; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field1_0_valid = out_carry_out_valid_R_1_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field1_0_bits_taskID = in_carry_in_R_1_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field1_0_bits_data = in_carry_in_R_1_data; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_InLiveOut_0_ready = ~ in_live_out_valid_R_0; // @[LoopBlock.scala 631:27]
  assign io_OutLiveOut_field0_0_valid = out_live_out_valid_R_0_0; // @[LoopBlock.scala 673:51]
  assign io_OutLiveOut_field0_0_bits_taskID = in_live_out_R_0_taskID; // @[LoopBlock.scala 672:50]
  assign io_OutLiveOut_field0_0_bits_data = in_live_out_R_0_data; // @[LoopBlock.scala 672:50]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
  assign _GEN_300 = _T_43 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_301 = _GEN_300 & _T_51; // @[LoopBlock.scala 932:19]
  assign _GEN_302 = _GEN_301 & _T_58; // @[LoopBlock.scala 932:19]
  assign _GEN_303 = _GEN_302 & loop_back_R_0_control; // @[LoopBlock.scala 932:19]
  assign _GEN_307 = loop_back_R_0_control == 1'h0; // @[LoopBlock.scala 950:19]
  assign _GEN_308 = _GEN_302 & _GEN_307; // @[LoopBlock.scala 950:19]
  assign _GEN_309 = _GEN_308 & loop_finish_R_0_control; // @[LoopBlock.scala 950:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_0_taskID = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_2_taskID = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_carry_in_R_1_taskID = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_carry_in_R_1_data = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_carry_in_valid_R_1 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_live_out_R_0_taskID = _RAND_23[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_live_out_R_0_data = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_live_out_valid_R_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  out_live_out_valid_R_0_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  out_live_out_fire_R_0_0 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  out_carry_out_valid_R_1_0 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_42[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  state = _RAND_46[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_43) begin
        if (_T_17) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_51) begin
          if (_T_17) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_17) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_17) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_17) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_51) begin
          if (_T_17) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_17) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_17) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_43) begin
        enable_valid_R <= _GEN_3;
      end else begin
        if (_T_51) begin
          enable_valid_R <= _GEN_3;
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_3;
            end
          end else begin
            enable_valid_R <= _GEN_3;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else begin
      if (_T_43) begin
        if (_T_19) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_19) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_19) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_19) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_19) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_19) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_19) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_19) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        loop_back_valid_R_0 <= _GEN_6;
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_21) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_21) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_21) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_21) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_7;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        loop_finish_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_43) begin
        if (_T_23) begin
          in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
        end
      end else begin
        if (_T_51) begin
          if (_T_23) begin
            in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_live_in_R_0_taskID <= 5'h0;
            end else begin
              if (_T_23) begin
                in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
              end
            end
          end else begin
            if (_T_23) begin
              in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_43) begin
        if (_T_23) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_51) begin
          if (_T_23) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_23) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_23) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_43) begin
        if (_T_25) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_51) begin
          if (_T_25) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_25) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_25) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_taskID <= 5'h0;
    end else begin
      if (_T_43) begin
        if (_T_27) begin
          in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
        end
      end else begin
        if (_T_51) begin
          if (_T_27) begin
            in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_live_in_R_2_taskID <= 5'h0;
            end else begin
              if (_T_27) begin
                in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
              end
            end
          end else begin
            if (_T_27) begin
              in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_43) begin
        if (_T_27) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_51) begin
          if (_T_27) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_27) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_27) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        in_live_in_valid_R_0 <= _GEN_13;
      end else begin
        if (_T_51) begin
          in_live_in_valid_R_0 <= _GEN_13;
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              in_live_in_valid_R_0 <= _GEN_13;
            end
          end else begin
            in_live_in_valid_R_0 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_43) begin
        in_live_in_valid_R_1 <= _GEN_17;
      end else begin
        if (_T_51) begin
          in_live_in_valid_R_1 <= _GEN_17;
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              in_live_in_valid_R_1 <= _GEN_17;
            end
          end else begin
            in_live_in_valid_R_1 <= _GEN_17;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_43) begin
        in_live_in_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_51) begin
          in_live_in_valid_R_2 <= _GEN_21;
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              in_live_in_valid_R_2 <= _GEN_21;
            end
          end else begin
            in_live_in_valid_R_2 <= _GEN_21;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_31) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_31) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_33) begin
        in_carry_in_R_1_taskID <= io_CarryDepenIn_1_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_1_data <= 32'h0;
    end else begin
      if (_T_33) begin
        in_carry_in_R_1_data <= io_CarryDepenIn_1_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        in_carry_in_valid_R_0 <= _GEN_29;
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_29;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_29;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_29;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_29;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_43) begin
        in_carry_in_valid_R_1 <= _GEN_33;
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_1 <= 1'h0;
            end else begin
              in_carry_in_valid_R_1 <= _GEN_33;
            end
          end else begin
            in_carry_in_valid_R_1 <= _GEN_33;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_carry_in_valid_R_1 <= 1'h0;
            end else begin
              in_carry_in_valid_R_1 <= _GEN_33;
            end
          end else begin
            in_carry_in_valid_R_1 <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      in_live_out_R_0_taskID <= 5'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          if (enable_R_control) begin
            if (_T_29) begin
              in_live_out_R_0_taskID <= io_InLiveOut_0_bits_taskID;
            end
          end else begin
            in_live_out_R_0_taskID <= 5'h0;
          end
        end else begin
          if (_T_29) begin
            in_live_out_R_0_taskID <= io_InLiveOut_0_bits_taskID;
          end
        end
      end else begin
        if (_T_29) begin
          in_live_out_R_0_taskID <= io_InLiveOut_0_bits_taskID;
        end
      end
    end
    if (reset) begin
      in_live_out_R_0_data <= 32'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          if (enable_R_control) begin
            if (_T_29) begin
              in_live_out_R_0_data <= io_InLiveOut_0_bits_data;
            end
          end else begin
            in_live_out_R_0_data <= 32'h0;
          end
        end else begin
          if (_T_29) begin
            in_live_out_R_0_data <= io_InLiveOut_0_bits_data;
          end
        end
      end else begin
        if (_T_29) begin
          in_live_out_R_0_data <= io_InLiveOut_0_bits_data;
        end
      end
    end
    if (reset) begin
      in_live_out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        in_live_out_valid_R_0 <= _GEN_25;
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              in_live_out_valid_R_0 <= 1'h0;
            end else begin
              in_live_out_valid_R_0 <= _GEN_25;
            end
          end else begin
            in_live_out_valid_R_0 <= _GEN_25;
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              in_live_out_valid_R_0 <= 1'h0;
            end else begin
              in_live_out_valid_R_0 <= _GEN_25;
            end
          end else begin
            in_live_out_valid_R_0 <= _GEN_25;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          out_live_in_valid_R_0_0 <= _GEN_50;
        end else begin
          if (_T_37) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            out_live_in_valid_R_0_0 <= _GEN_108;
          end else begin
            if (_T_37) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_37) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          out_live_in_valid_R_1_0 <= _GEN_51;
        end else begin
          if (_T_38) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            out_live_in_valid_R_1_0 <= _GEN_109;
          end else begin
            if (_T_38) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_38) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          out_live_in_valid_R_2_0 <= _GEN_52;
        end else begin
          if (_T_39) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            out_live_in_valid_R_2_0 <= _GEN_110;
          end else begin
            if (_T_39) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_39) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        out_live_in_fire_R_0_0 <= _GEN_39;
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_0 <= _GEN_39;
            end
          end else begin
            out_live_in_fire_R_0_0 <= _GEN_39;
          end
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_39;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        out_live_in_fire_R_1_0 <= _GEN_41;
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_0 <= _GEN_41;
            end
          end else begin
            out_live_in_fire_R_1_0 <= _GEN_41;
          end
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_41;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        out_live_in_fire_R_2_0 <= _GEN_43;
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_2_0 <= _GEN_43;
            end
          end else begin
            out_live_in_fire_R_2_0 <= _GEN_43;
          end
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_43;
        end
      end
    end
    if (reset) begin
      out_live_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          if (enable_R_control) begin
            if (_T_40) begin
              out_live_out_valid_R_0_0 <= 1'h0;
            end
          end else begin
            out_live_out_valid_R_0_0 <= 1'h1;
          end
        end else begin
          if (_T_40) begin
            out_live_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              if (_T_40) begin
                out_live_out_valid_R_0_0 <= 1'h0;
              end
            end else begin
              out_live_out_valid_R_0_0 <= _GEN_88;
            end
          end else begin
            if (_T_40) begin
              out_live_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_live_out_valid_R_0_0 <= _GEN_44;
        end
      end
    end
    if (reset) begin
      out_live_out_fire_R_0_0 <= 1'h0;
    end else begin
      out_live_out_fire_R_0_0 <= _GEN_45;
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          out_carry_out_valid_R_0_0 <= _GEN_53;
        end else begin
          if (_T_41) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            out_carry_out_valid_R_0_0 <= _GEN_111;
          end else begin
            if (_T_41) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_41) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          out_carry_out_valid_R_1_0 <= _GEN_54;
        end else begin
          if (_T_42) begin
            out_carry_out_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            out_carry_out_valid_R_1_0 <= _GEN_112;
          end else begin
            if (_T_42) begin
              out_carry_out_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_42) begin
            out_carry_out_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          active_loop_start_R_control <= _GEN_55;
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          active_loop_start_valid_R <= _GEN_57;
        end else begin
          if (_T_34) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            active_loop_start_valid_R <= _GEN_99;
          end else begin
            if (_T_34) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_34) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            active_loop_back_R_control <= _GEN_100;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          active_loop_back_valid_R <= _GEN_60;
        end else begin
          if (_T_35) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            active_loop_back_valid_R <= _GEN_102;
          end else begin
            if (_T_35) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_35) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 5'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          loop_exit_R_0_control <= _GEN_66;
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (!(loop_back_R_0_control)) begin
              loop_exit_R_0_control <= _GEN_94;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          if (enable_R_control) begin
            if (_T_36) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_36) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              if (_T_36) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              loop_exit_valid_R_0 <= _GEN_89;
            end
          end else begin
            if (_T_36) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_36;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_37;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_43) begin
        if (_T_46) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_51) begin
          if (_T_58) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_75) begin
            if (_T_76) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_303 & _T_65) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_0: Restarted fired @ %d\n",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 932:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_309 & _T_65) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_0: Output fired @ %d ",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 950:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_309 & _T_65) begin
          $fwrite(32'h80000002," Out[%d]: %d",1'h0,in_live_out_R_0_data); // @[LoopBlock.scala 953:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_309 & _T_65) begin
          $fwrite(32'h80000002,"\n"); // @[LoopBlock.scala 955:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [4:0]  io_InLiveIn_1_bits_taskID,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [31:0] io_InLiveIn_3_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [4:0]  io_OutLiveIn_field1_0_bits_taskID,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  output        io_CarryDepenIn_1_ready,
  input         io_CarryDepenIn_1_valid,
  input  [4:0]  io_CarryDepenIn_1_bits_taskID,
  input  [31:0] io_CarryDepenIn_1_bits_data,
  input         io_CarryDepenOut_field1_0_ready,
  output        io_CarryDepenOut_field1_0_valid,
  output [4:0]  io_CarryDepenOut_field1_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field1_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  output        io_InLiveOut_0_ready,
  input         io_InLiveOut_0_valid,
  input  [4:0]  io_InLiveOut_0_bits_taskID,
  input  [31:0] io_InLiveOut_0_bits_data,
  input         io_OutLiveOut_field0_0_ready,
  output        io_OutLiveOut_field0_0_valid,
  output [4:0]  io_OutLiveOut_field0_0_bits_taskID,
  output [31:0] io_OutLiveOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_2;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_3;
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_5;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_6;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_7;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_8;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [4:0] in_live_in_R_1_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_14;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_15;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_16;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_17;
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_18;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_19;
  reg [4:0] in_carry_in_R_1_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_20;
  reg [31:0] in_carry_in_R_1_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_21;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_22;
  reg  in_carry_in_valid_R_1; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_23;
  reg [4:0] in_live_out_R_0_taskID; // @[LoopBlock.scala 543:55]
  reg [31:0] _RAND_24;
  reg [31:0] in_live_out_R_0_data; // @[LoopBlock.scala 543:55]
  reg [31:0] _RAND_25;
  reg  in_live_out_valid_R_0; // @[LoopBlock.scala 544:61]
  reg [31:0] _RAND_26;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_27;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_28;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_29;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_30;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_31;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_32;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_33;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_34;
  reg  out_live_out_valid_R_0_0; // @[LoopBlock.scala 563:47]
  reg [31:0] _RAND_35;
  reg  out_live_out_fire_R_0_0; // @[LoopBlock.scala 567:47]
  reg [31:0] _RAND_36;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_37;
  reg  out_carry_out_valid_R_1_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_38;
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_39;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_40;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_41;
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_42;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_43;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_44;
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_45;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_46;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_47;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_48;
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[LoopBlock.scala 603:33]
  wire [4:0] _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_22; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_24; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_26; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_28; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_32; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[LoopBlock.scala 632:34]
  wire  _T_34; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[LoopBlock.scala 641:37]
  wire  _T_36; // @[Decoupled.scala 40:37]
  wire  _GEN_37; // @[LoopBlock.scala 641:37]
  wire  _T_37; // @[Decoupled.scala 40:37]
  wire  _GEN_38; // @[LoopBlock.scala 704:39]
  wire  _T_38; // @[Decoupled.scala 40:37]
  wire  _GEN_39; // @[LoopBlock.scala 708:38]
  wire  _T_39; // @[Decoupled.scala 40:37]
  wire  _GEN_40; // @[LoopBlock.scala 713:33]
  wire  _GEN_41; // @[LoopBlock.scala 713:33]
  wire  _T_40; // @[Decoupled.scala 40:37]
  wire  _GEN_42; // @[LoopBlock.scala 722:57]
  wire  _GEN_43; // @[LoopBlock.scala 722:57]
  wire  _T_41; // @[Decoupled.scala 40:37]
  wire  _GEN_44; // @[LoopBlock.scala 722:57]
  wire  _GEN_45; // @[LoopBlock.scala 722:57]
  wire  _T_42; // @[Decoupled.scala 40:37]
  wire  _GEN_46; // @[LoopBlock.scala 722:57]
  wire  _GEN_47; // @[LoopBlock.scala 722:57]
  wire  _T_43; // @[Decoupled.scala 40:37]
  wire  _GEN_48; // @[LoopBlock.scala 722:57]
  wire  _GEN_49; // @[LoopBlock.scala 722:57]
  wire  _T_44; // @[Decoupled.scala 40:37]
  wire  _GEN_50; // @[LoopBlock.scala 732:58]
  wire  _GEN_51; // @[LoopBlock.scala 732:58]
  wire  _T_45; // @[Decoupled.scala 40:37]
  wire  _GEN_52; // @[LoopBlock.scala 742:61]
  wire  _T_46; // @[Decoupled.scala 40:37]
  wire  _GEN_54; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_49;
  wire  _T_47; // @[Conditional.scala 37:30]
  wire  _T_48; // @[LoopBlock.scala 765:35]
  wire  _T_49; // @[LoopBlock.scala 765:35]
  wire  _T_50; // @[LoopBlock.scala 765:35]
  wire  _T_51; // @[LoopBlock.scala 869:28]
  wire  _GEN_56; // @[LoopBlock.scala 870:26]
  wire  _GEN_57; // @[LoopBlock.scala 870:26]
  wire  _GEN_58; // @[LoopBlock.scala 870:26]
  wire  _GEN_59; // @[LoopBlock.scala 870:26]
  wire  _GEN_60; // @[LoopBlock.scala 870:26]
  wire  _GEN_61; // @[LoopBlock.scala 870:26]
  wire  _GEN_62; // @[LoopBlock.scala 870:26]
  wire  _GEN_64; // @[LoopBlock.scala 870:26]
  wire  _GEN_67; // @[LoopBlock.scala 870:26]
  wire  _GEN_73; // @[LoopBlock.scala 870:26]
  wire  _T_56; // @[Conditional.scala 37:30]
  wire  _T_57; // @[LoopBlock.scala 898:30]
  wire  _T_58; // @[LoopBlock.scala 899:9]
  wire  _T_59; // @[LoopBlock.scala 828:26]
  wire  _T_60; // @[LoopBlock.scala 828:26]
  wire  _T_61; // @[LoopBlock.scala 828:26]
  wire  _T_62; // @[LoopBlock.scala 899:29]
  wire  _T_63; // @[LoopBlock.scala 783:40]
  wire  _T_64; // @[LoopBlock.scala 900:9]
  wire  _T_70; // @[LoopBlock.scala 932:19]
  wire  _T_71; // @[LoopBlock.scala 932:19]
  wire  _GEN_96; // @[LoopBlock.scala 936:64]
  wire  _GEN_97; // @[LoopBlock.scala 936:64]
  wire  _GEN_100; // @[LoopBlock.scala 936:64]
  wire  _GEN_102; // @[LoopBlock.scala 936:64]
  wire  _GEN_107; // @[LoopBlock.scala 903:56]
  wire  _GEN_108; // @[LoopBlock.scala 903:56]
  wire  _GEN_110; // @[LoopBlock.scala 903:56]
  wire  _GEN_117; // @[LoopBlock.scala 903:56]
  wire  _GEN_118; // @[LoopBlock.scala 903:56]
  wire  _GEN_119; // @[LoopBlock.scala 903:56]
  wire  _GEN_120; // @[LoopBlock.scala 903:56]
  wire  _GEN_121; // @[LoopBlock.scala 903:56]
  wire  _GEN_122; // @[LoopBlock.scala 903:56]
  wire  _T_81; // @[Conditional.scala 37:30]
  wire  _T_82; // @[LoopBlock.scala 963:27]
  wire  _GEN_332; // @[LoopBlock.scala 932:19]
  wire  _GEN_333; // @[LoopBlock.scala 932:19]
  wire  _GEN_334; // @[LoopBlock.scala 932:19]
  wire  _GEN_335; // @[LoopBlock.scala 932:19]
  wire  _GEN_339; // @[LoopBlock.scala 950:19]
  wire  _GEN_340; // @[LoopBlock.scala 950:19]
  wire  _GEN_341; // @[LoopBlock.scala 950:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_18 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_18 | enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_20 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_20 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_20 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_20 | loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_22 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_22 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_22 | loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_24 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_24 | in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_26 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_26 | in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_28 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_28 | in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_30 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_30 | in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_32 = io_InLiveOut_0_ready & io_InLiveOut_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_32 | in_live_out_valid_R_0; // @[LoopBlock.scala 632:34]
  assign _T_34 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_34 | in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_36 = io_CarryDepenIn_1_ready & io_CarryDepenIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_37 = _T_36 | in_carry_in_valid_R_1; // @[LoopBlock.scala 641:37]
  assign _T_37 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  assign _GEN_38 = _T_37 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_38 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  assign _GEN_39 = _T_38 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_39 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_40 = _T_39 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_41 = _T_39 | loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_40 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_42 = _T_40 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_43 = _T_40 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_41 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_44 = _T_41 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_45 = _T_41 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_42 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_46 = _T_42 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_47 = _T_42 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_43 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_48 = _T_43 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_49 = _T_43 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_44 = io_OutLiveOut_field0_0_ready & io_OutLiveOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_50 = _T_44 ? 1'h0 : out_live_out_valid_R_0_0; // @[LoopBlock.scala 732:58]
  assign _GEN_51 = _T_44 | out_live_out_fire_R_0_0; // @[LoopBlock.scala 732:58]
  assign _T_45 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_52 = _T_45 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_46 = io_CarryDepenOut_field1_0_ready & io_CarryDepenOut_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_54 = _T_46 ? 1'h0 : out_carry_out_valid_R_1_0; // @[LoopBlock.scala 742:61]
  assign _T_47 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_48 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_49 = _T_48 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_50 = _T_49 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_51 = _T_50 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_56 = enable_R_control | _GEN_42; // @[LoopBlock.scala 870:26]
  assign _GEN_57 = enable_R_control | _GEN_44; // @[LoopBlock.scala 870:26]
  assign _GEN_58 = enable_R_control | _GEN_46; // @[LoopBlock.scala 870:26]
  assign _GEN_59 = enable_R_control | _GEN_48; // @[LoopBlock.scala 870:26]
  assign _GEN_60 = enable_R_control | _GEN_52; // @[LoopBlock.scala 870:26]
  assign _GEN_61 = enable_R_control | _GEN_54; // @[LoopBlock.scala 870:26]
  assign _GEN_62 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_64 = enable_R_control | _GEN_38; // @[LoopBlock.scala 870:26]
  assign _GEN_67 = enable_R_control | _GEN_39; // @[LoopBlock.scala 870:26]
  assign _GEN_73 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 870:26]
  assign _T_56 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_57 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_58 = _T_57 & in_live_out_valid_R_0; // @[LoopBlock.scala 899:9]
  assign _T_59 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_60 = _T_59 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_61 = _T_60 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_62 = _T_58 & _T_61; // @[LoopBlock.scala 899:29]
  assign _T_63 = in_carry_in_valid_R_0 & in_carry_in_valid_R_1; // @[LoopBlock.scala 783:40]
  assign _T_64 = _T_62 & _T_63; // @[LoopBlock.scala 900:9]
  assign _T_70 = $unsigned(reset); // @[LoopBlock.scala 932:19]
  assign _T_71 = _T_70 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_96 = loop_finish_R_0_control | _GEN_50; // @[LoopBlock.scala 936:64]
  assign _GEN_97 = loop_finish_R_0_control | _GEN_40; // @[LoopBlock.scala 936:64]
  assign _GEN_100 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_102 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_107 = loop_back_R_0_control | _GEN_38; // @[LoopBlock.scala 903:56]
  assign _GEN_108 = loop_back_R_0_control | _GEN_100; // @[LoopBlock.scala 903:56]
  assign _GEN_110 = loop_back_R_0_control | _GEN_39; // @[LoopBlock.scala 903:56]
  assign _GEN_117 = loop_back_R_0_control | _GEN_42; // @[LoopBlock.scala 903:56]
  assign _GEN_118 = loop_back_R_0_control | _GEN_44; // @[LoopBlock.scala 903:56]
  assign _GEN_119 = loop_back_R_0_control | _GEN_46; // @[LoopBlock.scala 903:56]
  assign _GEN_120 = loop_back_R_0_control | _GEN_48; // @[LoopBlock.scala 903:56]
  assign _GEN_121 = loop_back_R_0_control | _GEN_52; // @[LoopBlock.scala 903:56]
  assign _GEN_122 = loop_back_R_0_control | _GEN_54; // @[LoopBlock.scala 903:56]
  assign _T_81 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_82 = loop_exit_fire_R_0 & out_live_out_fire_R_0_0; // @[LoopBlock.scala 963:27]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_taskID = in_live_in_R_1_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenIn_1_ready = ~ in_carry_in_valid_R_1; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field1_0_valid = out_carry_out_valid_R_1_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field1_0_bits_taskID = in_carry_in_R_1_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field1_0_bits_data = in_carry_in_R_1_data; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_InLiveOut_0_ready = ~ in_live_out_valid_R_0; // @[LoopBlock.scala 631:27]
  assign io_OutLiveOut_field0_0_valid = out_live_out_valid_R_0_0; // @[LoopBlock.scala 673:51]
  assign io_OutLiveOut_field0_0_bits_taskID = in_live_out_R_0_taskID; // @[LoopBlock.scala 672:50]
  assign io_OutLiveOut_field0_0_bits_data = in_live_out_R_0_data; // @[LoopBlock.scala 672:50]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
  assign _GEN_332 = _T_47 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_333 = _GEN_332 & _T_56; // @[LoopBlock.scala 932:19]
  assign _GEN_334 = _GEN_333 & _T_64; // @[LoopBlock.scala 932:19]
  assign _GEN_335 = _GEN_334 & loop_back_R_0_control; // @[LoopBlock.scala 932:19]
  assign _GEN_339 = loop_back_R_0_control == 1'h0; // @[LoopBlock.scala 950:19]
  assign _GEN_340 = _GEN_334 & _GEN_339; // @[LoopBlock.scala 950:19]
  assign _GEN_341 = _GEN_340 & loop_finish_R_0_control; // @[LoopBlock.scala 950:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_carry_in_R_1_taskID = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_carry_in_R_1_data = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_carry_in_valid_R_1 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_live_out_R_0_taskID = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_live_out_R_0_data = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  in_live_out_valid_R_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  out_live_out_valid_R_0_0 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  out_live_out_fire_R_0_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  out_carry_out_valid_R_1_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_39[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_42[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_45[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  state = _RAND_49[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_47) begin
        if (_T_18) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_56) begin
          if (_T_18) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_18) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_18) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_18) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_56) begin
          if (_T_18) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_18) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_18) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_47) begin
        enable_valid_R <= _GEN_3;
      end else begin
        if (_T_56) begin
          enable_valid_R <= _GEN_3;
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_3;
            end
          end else begin
            enable_valid_R <= _GEN_3;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else begin
      if (_T_47) begin
        if (_T_20) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_20) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_20) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_20) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_20) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_20) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_20) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_20) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        loop_back_valid_R_0 <= _GEN_6;
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_22) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_22) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_22) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_22) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_7;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        loop_finish_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_47) begin
        if (_T_24) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_56) begin
          if (_T_24) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_24) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_24) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_47) begin
        if (_T_26) begin
          in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
        end
      end else begin
        if (_T_56) begin
          if (_T_26) begin
            in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_in_R_1_taskID <= 5'h0;
            end else begin
              if (_T_26) begin
                in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
              end
            end
          end else begin
            if (_T_26) begin
              in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_47) begin
        if (_T_26) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_56) begin
          if (_T_26) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_26) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_26) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_47) begin
        if (_T_28) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_56) begin
          if (_T_28) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_28) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_28) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_47) begin
        if (_T_30) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_56) begin
          if (_T_30) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_30) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_30) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        in_live_in_valid_R_0 <= _GEN_13;
      end else begin
        if (_T_56) begin
          in_live_in_valid_R_0 <= _GEN_13;
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              in_live_in_valid_R_0 <= _GEN_13;
            end
          end else begin
            in_live_in_valid_R_0 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_47) begin
        in_live_in_valid_R_1 <= _GEN_17;
      end else begin
        if (_T_56) begin
          in_live_in_valid_R_1 <= _GEN_17;
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              in_live_in_valid_R_1 <= _GEN_17;
            end
          end else begin
            in_live_in_valid_R_1 <= _GEN_17;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_47) begin
        in_live_in_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_56) begin
          in_live_in_valid_R_2 <= _GEN_21;
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              in_live_in_valid_R_2 <= _GEN_21;
            end
          end else begin
            in_live_in_valid_R_2 <= _GEN_21;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_47) begin
        in_live_in_valid_R_3 <= _GEN_25;
      end else begin
        if (_T_56) begin
          in_live_in_valid_R_3 <= _GEN_25;
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              in_live_in_valid_R_3 <= _GEN_25;
            end
          end else begin
            in_live_in_valid_R_3 <= _GEN_25;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_34) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_34) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_36) begin
        in_carry_in_R_1_taskID <= io_CarryDepenIn_1_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_1_data <= 32'h0;
    end else begin
      if (_T_36) begin
        in_carry_in_R_1_data <= io_CarryDepenIn_1_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        in_carry_in_valid_R_0 <= _GEN_33;
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_33;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_33;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_33;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_47) begin
        in_carry_in_valid_R_1 <= _GEN_37;
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_1 <= 1'h0;
            end else begin
              in_carry_in_valid_R_1 <= _GEN_37;
            end
          end else begin
            in_carry_in_valid_R_1 <= _GEN_37;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_carry_in_valid_R_1 <= 1'h0;
            end else begin
              in_carry_in_valid_R_1 <= _GEN_37;
            end
          end else begin
            in_carry_in_valid_R_1 <= _GEN_37;
          end
        end
      end
    end
    if (reset) begin
      in_live_out_R_0_taskID <= 5'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          if (enable_R_control) begin
            if (_T_32) begin
              in_live_out_R_0_taskID <= io_InLiveOut_0_bits_taskID;
            end
          end else begin
            in_live_out_R_0_taskID <= 5'h0;
          end
        end else begin
          if (_T_32) begin
            in_live_out_R_0_taskID <= io_InLiveOut_0_bits_taskID;
          end
        end
      end else begin
        if (_T_32) begin
          in_live_out_R_0_taskID <= io_InLiveOut_0_bits_taskID;
        end
      end
    end
    if (reset) begin
      in_live_out_R_0_data <= 32'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          if (enable_R_control) begin
            if (_T_32) begin
              in_live_out_R_0_data <= io_InLiveOut_0_bits_data;
            end
          end else begin
            in_live_out_R_0_data <= 32'h0;
          end
        end else begin
          if (_T_32) begin
            in_live_out_R_0_data <= io_InLiveOut_0_bits_data;
          end
        end
      end else begin
        if (_T_32) begin
          in_live_out_R_0_data <= io_InLiveOut_0_bits_data;
        end
      end
    end
    if (reset) begin
      in_live_out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        in_live_out_valid_R_0 <= _GEN_29;
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              in_live_out_valid_R_0 <= 1'h0;
            end else begin
              in_live_out_valid_R_0 <= _GEN_29;
            end
          end else begin
            in_live_out_valid_R_0 <= _GEN_29;
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              in_live_out_valid_R_0 <= 1'h0;
            end else begin
              in_live_out_valid_R_0 <= _GEN_29;
            end
          end else begin
            in_live_out_valid_R_0 <= _GEN_29;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          out_live_in_valid_R_0_0 <= _GEN_56;
        end else begin
          if (_T_40) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            out_live_in_valid_R_0_0 <= _GEN_117;
          end else begin
            if (_T_40) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_40) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          out_live_in_valid_R_1_0 <= _GEN_57;
        end else begin
          if (_T_41) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            out_live_in_valid_R_1_0 <= _GEN_118;
          end else begin
            if (_T_41) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_41) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          out_live_in_valid_R_2_0 <= _GEN_58;
        end else begin
          if (_T_42) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            out_live_in_valid_R_2_0 <= _GEN_119;
          end else begin
            if (_T_42) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_42) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          out_live_in_valid_R_3_0 <= _GEN_59;
        end else begin
          if (_T_43) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            out_live_in_valid_R_3_0 <= _GEN_120;
          end else begin
            if (_T_43) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_43) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        out_live_in_fire_R_0_0 <= _GEN_43;
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_0 <= _GEN_43;
            end
          end else begin
            out_live_in_fire_R_0_0 <= _GEN_43;
          end
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_43;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        out_live_in_fire_R_1_0 <= _GEN_45;
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_0 <= _GEN_45;
            end
          end else begin
            out_live_in_fire_R_1_0 <= _GEN_45;
          end
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_45;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        out_live_in_fire_R_2_0 <= _GEN_47;
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_2_0 <= _GEN_47;
            end
          end else begin
            out_live_in_fire_R_2_0 <= _GEN_47;
          end
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_47;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        out_live_in_fire_R_3_0 <= _GEN_49;
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_3_0 <= _GEN_49;
            end
          end else begin
            out_live_in_fire_R_3_0 <= _GEN_49;
          end
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_49;
        end
      end
    end
    if (reset) begin
      out_live_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          if (enable_R_control) begin
            if (_T_44) begin
              out_live_out_valid_R_0_0 <= 1'h0;
            end
          end else begin
            out_live_out_valid_R_0_0 <= 1'h1;
          end
        end else begin
          if (_T_44) begin
            out_live_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              if (_T_44) begin
                out_live_out_valid_R_0_0 <= 1'h0;
              end
            end else begin
              out_live_out_valid_R_0_0 <= _GEN_96;
            end
          end else begin
            if (_T_44) begin
              out_live_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          out_live_out_valid_R_0_0 <= _GEN_50;
        end
      end
    end
    if (reset) begin
      out_live_out_fire_R_0_0 <= 1'h0;
    end else begin
      out_live_out_fire_R_0_0 <= _GEN_51;
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          out_carry_out_valid_R_0_0 <= _GEN_60;
        end else begin
          if (_T_45) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            out_carry_out_valid_R_0_0 <= _GEN_121;
          end else begin
            if (_T_45) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_45) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          out_carry_out_valid_R_1_0 <= _GEN_61;
        end else begin
          if (_T_46) begin
            out_carry_out_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            out_carry_out_valid_R_1_0 <= _GEN_122;
          end else begin
            if (_T_46) begin
              out_carry_out_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_46) begin
            out_carry_out_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          active_loop_start_R_control <= _GEN_62;
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          active_loop_start_valid_R <= _GEN_64;
        end else begin
          if (_T_37) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            active_loop_start_valid_R <= _GEN_107;
          end else begin
            if (_T_37) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_37) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            active_loop_back_R_control <= _GEN_108;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          active_loop_back_valid_R <= _GEN_67;
        end else begin
          if (_T_38) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            active_loop_back_valid_R <= _GEN_110;
          end else begin
            if (_T_38) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_38) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 5'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          loop_exit_R_0_control <= _GEN_73;
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (!(loop_back_R_0_control)) begin
              loop_exit_R_0_control <= _GEN_102;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          if (enable_R_control) begin
            if (_T_39) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_39) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              if (_T_39) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              loop_exit_valid_R_0 <= _GEN_97;
            end
          end else begin
            if (_T_39) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_40;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_41;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_47) begin
        if (_T_51) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_56) begin
          if (_T_64) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_81) begin
            if (_T_82) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_335 & _T_71) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_1: Restarted fired @ %d\n",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 932:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_341 & _T_71) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_1: Output fired @ %d ",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 950:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_341 & _T_71) begin
          $fwrite(32'h80000002," Out[%d]: %d",1'h0,in_live_out_R_0_data); // @[LoopBlock.scala 953:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_341 & _T_71) begin
          $fwrite(32'h80000002,"\n"); // @[LoopBlock.scala 955:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input         io_InLiveIn_1_bits_predicate,
  input  [4:0]  io_InLiveIn_1_bits_taskID,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [31:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [4:0]  io_InLiveIn_4_bits_taskID,
  input  [31:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input  [31:0] io_InLiveIn_5_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output [31:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [4:0]  io_OutLiveIn_field4_0_bits_taskID,
  output [31:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output        io_OutLiveIn_field1_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field1_0_bits_taskID,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field1_1_ready,
  output        io_OutLiveIn_field1_1_valid,
  output [4:0]  io_OutLiveIn_field1_1_bits_taskID,
  output [31:0] io_OutLiveIn_field1_1_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_2;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_3;
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_5;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_6;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_7;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_8;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg  in_live_in_R_1_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [4:0] in_live_in_R_1_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg [4:0] in_live_in_R_4_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_15;
  reg [31:0] in_live_in_R_4_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_16;
  reg [31:0] in_live_in_R_5_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_17;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_18;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_19;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_20;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_21;
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_22;
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_23;
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_24;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_25;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_26;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_27;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_28;
  reg  out_live_in_valid_R_1_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_29;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_30;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_31;
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_32;
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_33;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_34;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_35;
  reg  out_live_in_fire_R_1_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_36;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_37;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_38;
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_39;
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_40;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_41;
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_42;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_43;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_44;
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_45;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_46;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_47;
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_48;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_49;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_50;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_51;
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[LoopBlock.scala 603:33]
  wire [4:0] _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_22; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_24; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_26; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_28; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_32; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[LoopBlock.scala 623:33]
  wire  _T_34; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[LoopBlock.scala 623:33]
  wire  _T_36; // @[Decoupled.scala 40:37]
  wire  _GEN_37; // @[LoopBlock.scala 641:37]
  wire  _T_37; // @[Decoupled.scala 40:37]
  wire  _GEN_38; // @[LoopBlock.scala 704:39]
  wire  _T_38; // @[Decoupled.scala 40:37]
  wire  _GEN_39; // @[LoopBlock.scala 708:38]
  wire  _T_39; // @[Decoupled.scala 40:37]
  wire  _GEN_40; // @[LoopBlock.scala 713:33]
  wire  _GEN_41; // @[LoopBlock.scala 713:33]
  wire  _T_40; // @[Decoupled.scala 40:37]
  wire  _GEN_42; // @[LoopBlock.scala 722:57]
  wire  _GEN_43; // @[LoopBlock.scala 722:57]
  wire  _T_41; // @[Decoupled.scala 40:37]
  wire  _GEN_44; // @[LoopBlock.scala 722:57]
  wire  _GEN_45; // @[LoopBlock.scala 722:57]
  wire  _T_42; // @[Decoupled.scala 40:37]
  wire  _GEN_46; // @[LoopBlock.scala 722:57]
  wire  _GEN_47; // @[LoopBlock.scala 722:57]
  wire  _T_43; // @[Decoupled.scala 40:37]
  wire  _GEN_48; // @[LoopBlock.scala 722:57]
  wire  _GEN_49; // @[LoopBlock.scala 722:57]
  wire  _T_44; // @[Decoupled.scala 40:37]
  wire  _GEN_50; // @[LoopBlock.scala 722:57]
  wire  _GEN_51; // @[LoopBlock.scala 722:57]
  wire  _T_45; // @[Decoupled.scala 40:37]
  wire  _GEN_52; // @[LoopBlock.scala 722:57]
  wire  _GEN_53; // @[LoopBlock.scala 722:57]
  wire  _T_46; // @[Decoupled.scala 40:37]
  wire  _GEN_54; // @[LoopBlock.scala 722:57]
  wire  _GEN_55; // @[LoopBlock.scala 722:57]
  wire  _T_47; // @[Decoupled.scala 40:37]
  wire  _GEN_56; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_52;
  wire  _T_48; // @[Conditional.scala 37:30]
  wire  _T_49; // @[LoopBlock.scala 765:35]
  wire  _T_50; // @[LoopBlock.scala 765:35]
  wire  _T_51; // @[LoopBlock.scala 765:35]
  wire  _T_52; // @[LoopBlock.scala 765:35]
  wire  _T_53; // @[LoopBlock.scala 765:35]
  wire  _T_54; // @[LoopBlock.scala 869:28]
  wire  _GEN_58; // @[LoopBlock.scala 870:26]
  wire  _GEN_59; // @[LoopBlock.scala 870:26]
  wire  _GEN_60; // @[LoopBlock.scala 870:26]
  wire  _GEN_61; // @[LoopBlock.scala 870:26]
  wire  _GEN_62; // @[LoopBlock.scala 870:26]
  wire  _GEN_63; // @[LoopBlock.scala 870:26]
  wire  _GEN_64; // @[LoopBlock.scala 870:26]
  wire  _GEN_65; // @[LoopBlock.scala 870:26]
  wire  _GEN_66; // @[LoopBlock.scala 870:26]
  wire  _GEN_68; // @[LoopBlock.scala 870:26]
  wire  _GEN_71; // @[LoopBlock.scala 870:26]
  wire  _GEN_73; // @[LoopBlock.scala 870:26]
  wire  _T_58; // @[Conditional.scala 37:30]
  wire  _T_59; // @[LoopBlock.scala 898:30]
  wire  _T_61; // @[LoopBlock.scala 825:65]
  wire  _T_62; // @[LoopBlock.scala 828:26]
  wire  _T_63; // @[LoopBlock.scala 828:26]
  wire  _T_64; // @[LoopBlock.scala 828:26]
  wire  _T_65; // @[LoopBlock.scala 828:26]
  wire  _T_66; // @[LoopBlock.scala 828:26]
  wire  _T_67; // @[LoopBlock.scala 899:29]
  wire  _T_74; // @[LoopBlock.scala 932:19]
  wire  _T_75; // @[LoopBlock.scala 932:19]
  wire  _GEN_94; // @[LoopBlock.scala 936:64]
  wire  _GEN_97; // @[LoopBlock.scala 936:64]
  wire  _GEN_99; // @[LoopBlock.scala 936:64]
  wire  _GEN_104; // @[LoopBlock.scala 903:56]
  wire  _GEN_105; // @[LoopBlock.scala 903:56]
  wire  _GEN_107; // @[LoopBlock.scala 903:56]
  wire  _GEN_116; // @[LoopBlock.scala 903:56]
  wire  _GEN_117; // @[LoopBlock.scala 903:56]
  wire  _GEN_118; // @[LoopBlock.scala 903:56]
  wire  _GEN_119; // @[LoopBlock.scala 903:56]
  wire  _GEN_120; // @[LoopBlock.scala 903:56]
  wire  _GEN_121; // @[LoopBlock.scala 903:56]
  wire  _GEN_122; // @[LoopBlock.scala 903:56]
  wire  _GEN_123; // @[LoopBlock.scala 903:56]
  wire  _T_83; // @[Conditional.scala 37:30]
  wire  _GEN_358; // @[LoopBlock.scala 932:19]
  wire  _GEN_359; // @[LoopBlock.scala 932:19]
  wire  _GEN_360; // @[LoopBlock.scala 932:19]
  wire  _GEN_361; // @[LoopBlock.scala 932:19]
  wire  _GEN_365; // @[LoopBlock.scala 950:19]
  wire  _GEN_366; // @[LoopBlock.scala 950:19]
  wire  _GEN_367; // @[LoopBlock.scala 950:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_18 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_18 | enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_20 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_20 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_20 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_20 | loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_22 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_22 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_22 | loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_24 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_24 | in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_26 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_26 | in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_28 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_28 | in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_30 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_30 | in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_32 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_32 | in_live_in_valid_R_4; // @[LoopBlock.scala 623:33]
  assign _T_34 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_34 | in_live_in_valid_R_5; // @[LoopBlock.scala 623:33]
  assign _T_36 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_37 = _T_36 | in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_37 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  assign _GEN_38 = _T_37 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_38 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  assign _GEN_39 = _T_38 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_39 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_40 = _T_39 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_41 = _T_39 | loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_40 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_42 = _T_40 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_43 = _T_40 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_41 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_44 = _T_41 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_45 = _T_41 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_42 = io_OutLiveIn_field1_1_ready & io_OutLiveIn_field1_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_46 = _T_42 ? 1'h0 : out_live_in_valid_R_1_1; // @[LoopBlock.scala 722:57]
  assign _GEN_47 = _T_42 | out_live_in_fire_R_1_1; // @[LoopBlock.scala 722:57]
  assign _T_43 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_48 = _T_43 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_49 = _T_43 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_44 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_50 = _T_44 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_51 = _T_44 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_45 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_52 = _T_45 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 722:57]
  assign _GEN_53 = _T_45 | out_live_in_fire_R_4_0; // @[LoopBlock.scala 722:57]
  assign _T_46 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_54 = _T_46 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 722:57]
  assign _GEN_55 = _T_46 | out_live_in_fire_R_5_0; // @[LoopBlock.scala 722:57]
  assign _T_47 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_56 = _T_47 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_48 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_49 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_50 = _T_49 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_51 = _T_50 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_52 = _T_51 & in_live_in_valid_R_4; // @[LoopBlock.scala 765:35]
  assign _T_53 = _T_52 & in_live_in_valid_R_5; // @[LoopBlock.scala 765:35]
  assign _T_54 = _T_53 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_58 = enable_R_control | _GEN_42; // @[LoopBlock.scala 870:26]
  assign _GEN_59 = enable_R_control | _GEN_44; // @[LoopBlock.scala 870:26]
  assign _GEN_60 = enable_R_control | _GEN_46; // @[LoopBlock.scala 870:26]
  assign _GEN_61 = enable_R_control | _GEN_48; // @[LoopBlock.scala 870:26]
  assign _GEN_62 = enable_R_control | _GEN_50; // @[LoopBlock.scala 870:26]
  assign _GEN_63 = enable_R_control | _GEN_52; // @[LoopBlock.scala 870:26]
  assign _GEN_64 = enable_R_control | _GEN_54; // @[LoopBlock.scala 870:26]
  assign _GEN_65 = enable_R_control | _GEN_56; // @[LoopBlock.scala 870:26]
  assign _GEN_66 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_68 = enable_R_control | _GEN_38; // @[LoopBlock.scala 870:26]
  assign _GEN_71 = enable_R_control | _GEN_39; // @[LoopBlock.scala 870:26]
  assign _GEN_73 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 870:26]
  assign _T_58 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_59 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_61 = out_live_in_fire_R_1_0 & out_live_in_fire_R_1_1; // @[LoopBlock.scala 825:65]
  assign _T_62 = out_live_in_fire_R_0_0 & _T_61; // @[LoopBlock.scala 828:26]
  assign _T_63 = _T_62 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_64 = _T_63 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_65 = _T_64 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 828:26]
  assign _T_66 = _T_65 & out_live_in_fire_R_5_0; // @[LoopBlock.scala 828:26]
  assign _T_67 = _T_59 & _T_66; // @[LoopBlock.scala 899:29]
  assign _T_74 = $unsigned(reset); // @[LoopBlock.scala 932:19]
  assign _T_75 = _T_74 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_94 = loop_finish_R_0_control | _GEN_40; // @[LoopBlock.scala 936:64]
  assign _GEN_97 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_99 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_104 = loop_back_R_0_control | _GEN_38; // @[LoopBlock.scala 903:56]
  assign _GEN_105 = loop_back_R_0_control | _GEN_97; // @[LoopBlock.scala 903:56]
  assign _GEN_107 = loop_back_R_0_control | _GEN_39; // @[LoopBlock.scala 903:56]
  assign _GEN_116 = loop_back_R_0_control | _GEN_42; // @[LoopBlock.scala 903:56]
  assign _GEN_117 = loop_back_R_0_control | _GEN_44; // @[LoopBlock.scala 903:56]
  assign _GEN_118 = loop_back_R_0_control | _GEN_46; // @[LoopBlock.scala 903:56]
  assign _GEN_119 = loop_back_R_0_control | _GEN_48; // @[LoopBlock.scala 903:56]
  assign _GEN_120 = loop_back_R_0_control | _GEN_50; // @[LoopBlock.scala 903:56]
  assign _GEN_121 = loop_back_R_0_control | _GEN_52; // @[LoopBlock.scala 903:56]
  assign _GEN_122 = loop_back_R_0_control | _GEN_54; // @[LoopBlock.scala 903:56]
  assign _GEN_123 = loop_back_R_0_control | _GEN_56; // @[LoopBlock.scala 903:56]
  assign _T_83 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_4_ready = ~ in_live_in_valid_R_4; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_5_ready = ~ in_live_in_valid_R_5; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_0_bits_taskID = in_live_in_R_4_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_predicate = in_live_in_R_1_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_bits_taskID = in_live_in_R_1_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_1_valid = out_live_in_valid_R_1_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_1_bits_taskID = in_live_in_R_1_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_1_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
  assign _GEN_358 = _T_48 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_359 = _GEN_358 & _T_58; // @[LoopBlock.scala 932:19]
  assign _GEN_360 = _GEN_359 & _T_67; // @[LoopBlock.scala 932:19]
  assign _GEN_361 = _GEN_360 & loop_back_R_0_control; // @[LoopBlock.scala 932:19]
  assign _GEN_365 = loop_back_R_0_control == 1'h0; // @[LoopBlock.scala 950:19]
  assign _GEN_366 = _GEN_360 & _GEN_365; // @[LoopBlock.scala 950:19]
  assign _GEN_367 = _GEN_366 & loop_finish_R_0_control; // @[LoopBlock.scala 950:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_predicate = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_1_taskID = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_R_4_taskID = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_R_4_data = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_R_5_data = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_live_in_valid_R_1_1 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  out_live_in_fire_R_1_1 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_42[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_45[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_48[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  state = _RAND_52[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_48) begin
        if (_T_18) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_58) begin
          if (_T_18) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_18) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_18) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_18) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_58) begin
          if (_T_18) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_18) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_18) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_48) begin
        enable_valid_R <= _GEN_3;
      end else begin
        if (_T_58) begin
          enable_valid_R <= _GEN_3;
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_3;
            end
          end else begin
            enable_valid_R <= _GEN_3;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else begin
      if (_T_48) begin
        if (_T_20) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_20) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_20) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_20) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_20) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_20) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_20) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_20) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        loop_back_valid_R_0 <= _GEN_6;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_22) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_22) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_22) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_22) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_7;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        loop_finish_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_48) begin
        if (_T_24) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_58) begin
          if (_T_24) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_24) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_24) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_predicate <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_26) begin
          in_live_in_R_1_predicate <= io_InLiveIn_1_bits_predicate;
        end
      end else begin
        if (_T_58) begin
          if (_T_26) begin
            in_live_in_R_1_predicate <= io_InLiveIn_1_bits_predicate;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_predicate <= 1'h0;
            end else begin
              if (_T_26) begin
                in_live_in_R_1_predicate <= io_InLiveIn_1_bits_predicate;
              end
            end
          end else begin
            if (_T_26) begin
              in_live_in_R_1_predicate <= io_InLiveIn_1_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_48) begin
        if (_T_26) begin
          in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
        end
      end else begin
        if (_T_58) begin
          if (_T_26) begin
            in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_taskID <= 5'h0;
            end else begin
              if (_T_26) begin
                in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
              end
            end
          end else begin
            if (_T_26) begin
              in_live_in_R_1_taskID <= io_InLiveIn_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_48) begin
        if (_T_26) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_58) begin
          if (_T_26) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_26) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_26) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_48) begin
        if (_T_28) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_58) begin
          if (_T_28) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_28) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_28) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_48) begin
        if (_T_30) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_58) begin
          if (_T_30) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_30) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_30) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_taskID <= 5'h0;
    end else begin
      if (_T_48) begin
        if (_T_32) begin
          in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
        end
      end else begin
        if (_T_58) begin
          if (_T_32) begin
            in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_taskID <= 5'h0;
            end else begin
              if (_T_32) begin
                in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
              end
            end
          end else begin
            if (_T_32) begin
              in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_data <= 32'h0;
    end else begin
      if (_T_48) begin
        if (_T_32) begin
          in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
        end
      end else begin
        if (_T_58) begin
          if (_T_32) begin
            in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_data <= 32'h0;
            end else begin
              if (_T_32) begin
                in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
              end
            end
          end else begin
            if (_T_32) begin
              in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_data <= 32'h0;
    end else begin
      if (_T_48) begin
        if (_T_34) begin
          in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
        end
      end else begin
        if (_T_58) begin
          if (_T_34) begin
            in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_data <= 32'h0;
            end else begin
              if (_T_34) begin
                in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
              end
            end
          end else begin
            if (_T_34) begin
              in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        in_live_in_valid_R_0 <= _GEN_13;
      end else begin
        if (_T_58) begin
          in_live_in_valid_R_0 <= _GEN_13;
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              in_live_in_valid_R_0 <= _GEN_13;
            end
          end else begin
            in_live_in_valid_R_0 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_48) begin
        in_live_in_valid_R_1 <= _GEN_17;
      end else begin
        if (_T_58) begin
          in_live_in_valid_R_1 <= _GEN_17;
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              in_live_in_valid_R_1 <= _GEN_17;
            end
          end else begin
            in_live_in_valid_R_1 <= _GEN_17;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_48) begin
        in_live_in_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_58) begin
          in_live_in_valid_R_2 <= _GEN_21;
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              in_live_in_valid_R_2 <= _GEN_21;
            end
          end else begin
            in_live_in_valid_R_2 <= _GEN_21;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_48) begin
        in_live_in_valid_R_3 <= _GEN_25;
      end else begin
        if (_T_58) begin
          in_live_in_valid_R_3 <= _GEN_25;
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              in_live_in_valid_R_3 <= _GEN_25;
            end
          end else begin
            in_live_in_valid_R_3 <= _GEN_25;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else begin
      if (_T_48) begin
        in_live_in_valid_R_4 <= _GEN_29;
      end else begin
        if (_T_58) begin
          in_live_in_valid_R_4 <= _GEN_29;
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_4 <= 1'h0;
            end else begin
              in_live_in_valid_R_4 <= _GEN_29;
            end
          end else begin
            in_live_in_valid_R_4 <= _GEN_29;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else begin
      if (_T_48) begin
        in_live_in_valid_R_5 <= _GEN_33;
      end else begin
        if (_T_58) begin
          in_live_in_valid_R_5 <= _GEN_33;
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_5 <= 1'h0;
            end else begin
              in_live_in_valid_R_5 <= _GEN_33;
            end
          end else begin
            in_live_in_valid_R_5 <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_36) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_36) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        in_carry_in_valid_R_0 <= _GEN_37;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_37;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_37;
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_37;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_37;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          out_live_in_valid_R_0_0 <= _GEN_58;
        end else begin
          if (_T_40) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            out_live_in_valid_R_0_0 <= _GEN_116;
          end else begin
            if (_T_40) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_40) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          out_live_in_valid_R_1_0 <= _GEN_59;
        end else begin
          if (_T_41) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            out_live_in_valid_R_1_0 <= _GEN_117;
          end else begin
            if (_T_41) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_41) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_1 <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          out_live_in_valid_R_1_1 <= _GEN_60;
        end else begin
          if (_T_42) begin
            out_live_in_valid_R_1_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            out_live_in_valid_R_1_1 <= _GEN_118;
          end else begin
            if (_T_42) begin
              out_live_in_valid_R_1_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_42) begin
            out_live_in_valid_R_1_1 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          out_live_in_valid_R_2_0 <= _GEN_61;
        end else begin
          if (_T_43) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            out_live_in_valid_R_2_0 <= _GEN_119;
          end else begin
            if (_T_43) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_43) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          out_live_in_valid_R_3_0 <= _GEN_62;
        end else begin
          if (_T_44) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            out_live_in_valid_R_3_0 <= _GEN_120;
          end else begin
            if (_T_44) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_44) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          out_live_in_valid_R_4_0 <= _GEN_63;
        end else begin
          if (_T_45) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            out_live_in_valid_R_4_0 <= _GEN_121;
          end else begin
            if (_T_45) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_45) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          out_live_in_valid_R_5_0 <= _GEN_64;
        end else begin
          if (_T_46) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            out_live_in_valid_R_5_0 <= _GEN_122;
          end else begin
            if (_T_46) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_46) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        out_live_in_fire_R_0_0 <= _GEN_43;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_0 <= _GEN_43;
            end
          end else begin
            out_live_in_fire_R_0_0 <= _GEN_43;
          end
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_43;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        out_live_in_fire_R_1_0 <= _GEN_45;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_0 <= _GEN_45;
            end
          end else begin
            out_live_in_fire_R_1_0 <= _GEN_45;
          end
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_45;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_1 <= 1'h0;
    end else begin
      if (_T_48) begin
        out_live_in_fire_R_1_1 <= _GEN_47;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_1 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_1 <= _GEN_47;
            end
          end else begin
            out_live_in_fire_R_1_1 <= _GEN_47;
          end
        end else begin
          out_live_in_fire_R_1_1 <= _GEN_47;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        out_live_in_fire_R_2_0 <= _GEN_49;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_2_0 <= _GEN_49;
            end
          end else begin
            out_live_in_fire_R_2_0 <= _GEN_49;
          end
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_49;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        out_live_in_fire_R_3_0 <= _GEN_51;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_3_0 <= _GEN_51;
            end
          end else begin
            out_live_in_fire_R_3_0 <= _GEN_51;
          end
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_51;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        out_live_in_fire_R_4_0 <= _GEN_53;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_4_0 <= _GEN_53;
            end
          end else begin
            out_live_in_fire_R_4_0 <= _GEN_53;
          end
        end else begin
          out_live_in_fire_R_4_0 <= _GEN_53;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        out_live_in_fire_R_5_0 <= _GEN_55;
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_5_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_5_0 <= _GEN_55;
            end
          end else begin
            out_live_in_fire_R_5_0 <= _GEN_55;
          end
        end else begin
          out_live_in_fire_R_5_0 <= _GEN_55;
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          out_carry_out_valid_R_0_0 <= _GEN_65;
        end else begin
          if (_T_47) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            out_carry_out_valid_R_0_0 <= _GEN_123;
          end else begin
            if (_T_47) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_47) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          active_loop_start_R_control <= _GEN_66;
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          active_loop_start_valid_R <= _GEN_68;
        end else begin
          if (_T_37) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            active_loop_start_valid_R <= _GEN_104;
          end else begin
            if (_T_37) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_37) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            active_loop_back_R_control <= _GEN_105;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          active_loop_back_valid_R <= _GEN_71;
        end else begin
          if (_T_38) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            active_loop_back_valid_R <= _GEN_107;
          end else begin
            if (_T_38) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_38) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 5'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          loop_exit_R_0_control <= _GEN_73;
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (!(loop_back_R_0_control)) begin
              loop_exit_R_0_control <= _GEN_99;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          if (enable_R_control) begin
            if (_T_39) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_39) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              if (_T_39) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              loop_exit_valid_R_0 <= _GEN_94;
            end
          end else begin
            if (_T_39) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_40;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_41;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_48) begin
        if (_T_54) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_58) begin
          if (_T_67) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_83) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_361 & _T_75) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_2: Restarted fired @ %d\n",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 932:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & _T_75) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_2: Output fired @ %d ",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 950:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_367 & _T_75) begin
          $fwrite(32'h80000002,"\n"); // @[LoopBlock.scala 955:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [31:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [4:0]  io_InLiveIn_4_bits_taskID,
  input  [31:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input  [4:0]  io_InLiveIn_5_bits_taskID,
  input  [31:0] io_InLiveIn_5_bits_data,
  output        io_InLiveIn_6_ready,
  input         io_InLiveIn_6_valid,
  input  [31:0] io_InLiveIn_6_bits_data,
  output        io_InLiveIn_7_ready,
  input         io_InLiveIn_7_valid,
  input  [31:0] io_InLiveIn_7_bits_data,
  output        io_InLiveIn_8_ready,
  input         io_InLiveIn_8_valid,
  input  [4:0]  io_InLiveIn_8_bits_taskID,
  input  [31:0] io_InLiveIn_8_bits_data,
  input         io_OutLiveIn_field8_0_ready,
  output        io_OutLiveIn_field8_0_valid,
  output [4:0]  io_OutLiveIn_field8_0_bits_taskID,
  output [31:0] io_OutLiveIn_field8_0_bits_data,
  input         io_OutLiveIn_field8_1_ready,
  output        io_OutLiveIn_field8_1_valid,
  output [31:0] io_OutLiveIn_field8_1_bits_data,
  input         io_OutLiveIn_field7_0_ready,
  output        io_OutLiveIn_field7_0_valid,
  output [31:0] io_OutLiveIn_field7_0_bits_data,
  input         io_OutLiveIn_field6_0_ready,
  output        io_OutLiveIn_field6_0_valid,
  output [31:0] io_OutLiveIn_field6_0_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output [4:0]  io_OutLiveIn_field5_0_bits_taskID,
  output [31:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [4:0]  io_OutLiveIn_field4_0_bits_taskID,
  output [31:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_2;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_3;
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_5;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_6;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_7;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_8;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [4:0] in_live_in_R_4_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [31:0] in_live_in_R_4_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg [4:0] in_live_in_R_5_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_15;
  reg [31:0] in_live_in_R_5_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_16;
  reg [31:0] in_live_in_R_6_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_17;
  reg [31:0] in_live_in_R_7_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_18;
  reg [4:0] in_live_in_R_8_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_19;
  reg [31:0] in_live_in_R_8_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_20;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_21;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_22;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_23;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_24;
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_25;
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_26;
  reg  in_live_in_valid_R_6; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_27;
  reg  in_live_in_valid_R_7; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_28;
  reg  in_live_in_valid_R_8; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_29;
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_30;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_31;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_32;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_33;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_34;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_35;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_36;
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_37;
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_38;
  reg  out_live_in_valid_R_6_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_39;
  reg  out_live_in_valid_R_7_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_40;
  reg  out_live_in_valid_R_8_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_41;
  reg  out_live_in_valid_R_8_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_42;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_43;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_44;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_45;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_46;
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_47;
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_48;
  reg  out_live_in_fire_R_6_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_49;
  reg  out_live_in_fire_R_7_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_50;
  reg  out_live_in_fire_R_8_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_51;
  reg  out_live_in_fire_R_8_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_52;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_53;
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_54;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_55;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_56;
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_57;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_58;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_59;
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_60;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_61;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_62;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_63;
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[LoopBlock.scala 603:33]
  wire [4:0] _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_25; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_27; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_29; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_31; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_33; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_35; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[LoopBlock.scala 623:33]
  wire  _T_37; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[LoopBlock.scala 623:33]
  wire  _T_39; // @[Decoupled.scala 40:37]
  wire  _GEN_37; // @[LoopBlock.scala 623:33]
  wire  _T_41; // @[Decoupled.scala 40:37]
  wire  _GEN_41; // @[LoopBlock.scala 623:33]
  wire  _T_43; // @[Decoupled.scala 40:37]
  wire  _GEN_45; // @[LoopBlock.scala 623:33]
  wire  _T_45; // @[Decoupled.scala 40:37]
  wire  _GEN_49; // @[LoopBlock.scala 641:37]
  wire  _T_46; // @[Decoupled.scala 40:37]
  wire  _GEN_50; // @[LoopBlock.scala 704:39]
  wire  _T_47; // @[Decoupled.scala 40:37]
  wire  _GEN_51; // @[LoopBlock.scala 708:38]
  wire  _T_48; // @[Decoupled.scala 40:37]
  wire  _GEN_52; // @[LoopBlock.scala 713:33]
  wire  _GEN_53; // @[LoopBlock.scala 713:33]
  wire  _T_49; // @[Decoupled.scala 40:37]
  wire  _GEN_54; // @[LoopBlock.scala 722:57]
  wire  _GEN_55; // @[LoopBlock.scala 722:57]
  wire  _T_50; // @[Decoupled.scala 40:37]
  wire  _GEN_56; // @[LoopBlock.scala 722:57]
  wire  _GEN_57; // @[LoopBlock.scala 722:57]
  wire  _T_51; // @[Decoupled.scala 40:37]
  wire  _GEN_58; // @[LoopBlock.scala 722:57]
  wire  _GEN_59; // @[LoopBlock.scala 722:57]
  wire  _T_52; // @[Decoupled.scala 40:37]
  wire  _GEN_60; // @[LoopBlock.scala 722:57]
  wire  _GEN_61; // @[LoopBlock.scala 722:57]
  wire  _T_53; // @[Decoupled.scala 40:37]
  wire  _GEN_62; // @[LoopBlock.scala 722:57]
  wire  _GEN_63; // @[LoopBlock.scala 722:57]
  wire  _T_54; // @[Decoupled.scala 40:37]
  wire  _GEN_64; // @[LoopBlock.scala 722:57]
  wire  _GEN_65; // @[LoopBlock.scala 722:57]
  wire  _T_55; // @[Decoupled.scala 40:37]
  wire  _GEN_66; // @[LoopBlock.scala 722:57]
  wire  _GEN_67; // @[LoopBlock.scala 722:57]
  wire  _T_56; // @[Decoupled.scala 40:37]
  wire  _GEN_68; // @[LoopBlock.scala 722:57]
  wire  _GEN_69; // @[LoopBlock.scala 722:57]
  wire  _T_57; // @[Decoupled.scala 40:37]
  wire  _GEN_70; // @[LoopBlock.scala 722:57]
  wire  _GEN_71; // @[LoopBlock.scala 722:57]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire  _GEN_72; // @[LoopBlock.scala 722:57]
  wire  _GEN_73; // @[LoopBlock.scala 722:57]
  wire  _T_59; // @[Decoupled.scala 40:37]
  wire  _GEN_74; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_64;
  wire  _T_60; // @[Conditional.scala 37:30]
  wire  _T_61; // @[LoopBlock.scala 765:35]
  wire  _T_62; // @[LoopBlock.scala 765:35]
  wire  _T_63; // @[LoopBlock.scala 765:35]
  wire  _T_64; // @[LoopBlock.scala 765:35]
  wire  _T_65; // @[LoopBlock.scala 765:35]
  wire  _T_66; // @[LoopBlock.scala 765:35]
  wire  _T_67; // @[LoopBlock.scala 765:35]
  wire  _T_68; // @[LoopBlock.scala 765:35]
  wire  _T_69; // @[LoopBlock.scala 869:28]
  wire  _GEN_76; // @[LoopBlock.scala 870:26]
  wire  _GEN_77; // @[LoopBlock.scala 870:26]
  wire  _GEN_78; // @[LoopBlock.scala 870:26]
  wire  _GEN_79; // @[LoopBlock.scala 870:26]
  wire  _GEN_80; // @[LoopBlock.scala 870:26]
  wire  _GEN_81; // @[LoopBlock.scala 870:26]
  wire  _GEN_82; // @[LoopBlock.scala 870:26]
  wire  _GEN_83; // @[LoopBlock.scala 870:26]
  wire  _GEN_84; // @[LoopBlock.scala 870:26]
  wire  _GEN_85; // @[LoopBlock.scala 870:26]
  wire  _GEN_86; // @[LoopBlock.scala 870:26]
  wire  _GEN_87; // @[LoopBlock.scala 870:26]
  wire  _GEN_89; // @[LoopBlock.scala 870:26]
  wire  _GEN_92; // @[LoopBlock.scala 870:26]
  wire  _GEN_94; // @[LoopBlock.scala 870:26]
  wire  _T_73; // @[Conditional.scala 37:30]
  wire  _T_74; // @[LoopBlock.scala 898:30]
  wire  _T_76; // @[LoopBlock.scala 825:65]
  wire  _T_77; // @[LoopBlock.scala 828:26]
  wire  _T_78; // @[LoopBlock.scala 828:26]
  wire  _T_79; // @[LoopBlock.scala 828:26]
  wire  _T_80; // @[LoopBlock.scala 828:26]
  wire  _T_81; // @[LoopBlock.scala 828:26]
  wire  _T_82; // @[LoopBlock.scala 828:26]
  wire  _T_83; // @[LoopBlock.scala 828:26]
  wire  _T_84; // @[LoopBlock.scala 828:26]
  wire  _T_85; // @[LoopBlock.scala 899:29]
  wire  _T_92; // @[LoopBlock.scala 932:19]
  wire  _T_93; // @[LoopBlock.scala 932:19]
  wire  _GEN_118; // @[LoopBlock.scala 936:64]
  wire  _GEN_121; // @[LoopBlock.scala 936:64]
  wire  _GEN_123; // @[LoopBlock.scala 936:64]
  wire  _GEN_128; // @[LoopBlock.scala 903:56]
  wire  _GEN_129; // @[LoopBlock.scala 903:56]
  wire  _GEN_131; // @[LoopBlock.scala 903:56]
  wire  _GEN_143; // @[LoopBlock.scala 903:56]
  wire  _GEN_144; // @[LoopBlock.scala 903:56]
  wire  _GEN_145; // @[LoopBlock.scala 903:56]
  wire  _GEN_146; // @[LoopBlock.scala 903:56]
  wire  _GEN_147; // @[LoopBlock.scala 903:56]
  wire  _GEN_148; // @[LoopBlock.scala 903:56]
  wire  _GEN_149; // @[LoopBlock.scala 903:56]
  wire  _GEN_150; // @[LoopBlock.scala 903:56]
  wire  _GEN_151; // @[LoopBlock.scala 903:56]
  wire  _GEN_152; // @[LoopBlock.scala 903:56]
  wire  _GEN_153; // @[LoopBlock.scala 903:56]
  wire  _T_101; // @[Conditional.scala 37:30]
  wire  _GEN_454; // @[LoopBlock.scala 932:19]
  wire  _GEN_455; // @[LoopBlock.scala 932:19]
  wire  _GEN_456; // @[LoopBlock.scala 932:19]
  wire  _GEN_457; // @[LoopBlock.scala 932:19]
  wire  _GEN_461; // @[LoopBlock.scala 950:19]
  wire  _GEN_462; // @[LoopBlock.scala 950:19]
  wire  _GEN_463; // @[LoopBlock.scala 950:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_21 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_21 | enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_23 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_23 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_23 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_23 | loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_25 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_25 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_25 | loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_27 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_27 | in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_29 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_29 | in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_31 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_31 | in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_33 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_33 | in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_35 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_35 | in_live_in_valid_R_4; // @[LoopBlock.scala 623:33]
  assign _T_37 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_37 | in_live_in_valid_R_5; // @[LoopBlock.scala 623:33]
  assign _T_39 = io_InLiveIn_6_ready & io_InLiveIn_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_37 = _T_39 | in_live_in_valid_R_6; // @[LoopBlock.scala 623:33]
  assign _T_41 = io_InLiveIn_7_ready & io_InLiveIn_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_41 = _T_41 | in_live_in_valid_R_7; // @[LoopBlock.scala 623:33]
  assign _T_43 = io_InLiveIn_8_ready & io_InLiveIn_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_45 = _T_43 | in_live_in_valid_R_8; // @[LoopBlock.scala 623:33]
  assign _T_45 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_49 = _T_45 | in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_46 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  assign _GEN_50 = _T_46 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_47 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  assign _GEN_51 = _T_47 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_48 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_52 = _T_48 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_53 = _T_48 | loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_49 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_54 = _T_49 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_55 = _T_49 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_50 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_56 = _T_50 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_57 = _T_50 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_51 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_58 = _T_51 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_59 = _T_51 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_52 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_60 = _T_52 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_61 = _T_52 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_53 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_62 = _T_53 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 722:57]
  assign _GEN_63 = _T_53 | out_live_in_fire_R_4_0; // @[LoopBlock.scala 722:57]
  assign _T_54 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_64 = _T_54 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 722:57]
  assign _GEN_65 = _T_54 | out_live_in_fire_R_5_0; // @[LoopBlock.scala 722:57]
  assign _T_55 = io_OutLiveIn_field6_0_ready & io_OutLiveIn_field6_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_66 = _T_55 ? 1'h0 : out_live_in_valid_R_6_0; // @[LoopBlock.scala 722:57]
  assign _GEN_67 = _T_55 | out_live_in_fire_R_6_0; // @[LoopBlock.scala 722:57]
  assign _T_56 = io_OutLiveIn_field7_0_ready & io_OutLiveIn_field7_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_68 = _T_56 ? 1'h0 : out_live_in_valid_R_7_0; // @[LoopBlock.scala 722:57]
  assign _GEN_69 = _T_56 | out_live_in_fire_R_7_0; // @[LoopBlock.scala 722:57]
  assign _T_57 = io_OutLiveIn_field8_0_ready & io_OutLiveIn_field8_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_70 = _T_57 ? 1'h0 : out_live_in_valid_R_8_0; // @[LoopBlock.scala 722:57]
  assign _GEN_71 = _T_57 | out_live_in_fire_R_8_0; // @[LoopBlock.scala 722:57]
  assign _T_58 = io_OutLiveIn_field8_1_ready & io_OutLiveIn_field8_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_72 = _T_58 ? 1'h0 : out_live_in_valid_R_8_1; // @[LoopBlock.scala 722:57]
  assign _GEN_73 = _T_58 | out_live_in_fire_R_8_1; // @[LoopBlock.scala 722:57]
  assign _T_59 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_74 = _T_59 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_60 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_61 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_62 = _T_61 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_63 = _T_62 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_64 = _T_63 & in_live_in_valid_R_4; // @[LoopBlock.scala 765:35]
  assign _T_65 = _T_64 & in_live_in_valid_R_5; // @[LoopBlock.scala 765:35]
  assign _T_66 = _T_65 & in_live_in_valid_R_6; // @[LoopBlock.scala 765:35]
  assign _T_67 = _T_66 & in_live_in_valid_R_7; // @[LoopBlock.scala 765:35]
  assign _T_68 = _T_67 & in_live_in_valid_R_8; // @[LoopBlock.scala 765:35]
  assign _T_69 = _T_68 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_76 = enable_R_control | _GEN_54; // @[LoopBlock.scala 870:26]
  assign _GEN_77 = enable_R_control | _GEN_56; // @[LoopBlock.scala 870:26]
  assign _GEN_78 = enable_R_control | _GEN_58; // @[LoopBlock.scala 870:26]
  assign _GEN_79 = enable_R_control | _GEN_60; // @[LoopBlock.scala 870:26]
  assign _GEN_80 = enable_R_control | _GEN_62; // @[LoopBlock.scala 870:26]
  assign _GEN_81 = enable_R_control | _GEN_64; // @[LoopBlock.scala 870:26]
  assign _GEN_82 = enable_R_control | _GEN_66; // @[LoopBlock.scala 870:26]
  assign _GEN_83 = enable_R_control | _GEN_68; // @[LoopBlock.scala 870:26]
  assign _GEN_84 = enable_R_control | _GEN_70; // @[LoopBlock.scala 870:26]
  assign _GEN_85 = enable_R_control | _GEN_72; // @[LoopBlock.scala 870:26]
  assign _GEN_86 = enable_R_control | _GEN_74; // @[LoopBlock.scala 870:26]
  assign _GEN_87 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_89 = enable_R_control | _GEN_50; // @[LoopBlock.scala 870:26]
  assign _GEN_92 = enable_R_control | _GEN_51; // @[LoopBlock.scala 870:26]
  assign _GEN_94 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 870:26]
  assign _T_73 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_74 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_76 = out_live_in_fire_R_8_0 & out_live_in_fire_R_8_1; // @[LoopBlock.scala 825:65]
  assign _T_77 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_78 = _T_77 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_79 = _T_78 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_80 = _T_79 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 828:26]
  assign _T_81 = _T_80 & out_live_in_fire_R_5_0; // @[LoopBlock.scala 828:26]
  assign _T_82 = _T_81 & out_live_in_fire_R_6_0; // @[LoopBlock.scala 828:26]
  assign _T_83 = _T_82 & out_live_in_fire_R_7_0; // @[LoopBlock.scala 828:26]
  assign _T_84 = _T_83 & _T_76; // @[LoopBlock.scala 828:26]
  assign _T_85 = _T_74 & _T_84; // @[LoopBlock.scala 899:29]
  assign _T_92 = $unsigned(reset); // @[LoopBlock.scala 932:19]
  assign _T_93 = _T_92 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_118 = loop_finish_R_0_control | _GEN_52; // @[LoopBlock.scala 936:64]
  assign _GEN_121 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_123 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_128 = loop_back_R_0_control | _GEN_50; // @[LoopBlock.scala 903:56]
  assign _GEN_129 = loop_back_R_0_control | _GEN_121; // @[LoopBlock.scala 903:56]
  assign _GEN_131 = loop_back_R_0_control | _GEN_51; // @[LoopBlock.scala 903:56]
  assign _GEN_143 = loop_back_R_0_control | _GEN_54; // @[LoopBlock.scala 903:56]
  assign _GEN_144 = loop_back_R_0_control | _GEN_56; // @[LoopBlock.scala 903:56]
  assign _GEN_145 = loop_back_R_0_control | _GEN_58; // @[LoopBlock.scala 903:56]
  assign _GEN_146 = loop_back_R_0_control | _GEN_60; // @[LoopBlock.scala 903:56]
  assign _GEN_147 = loop_back_R_0_control | _GEN_62; // @[LoopBlock.scala 903:56]
  assign _GEN_148 = loop_back_R_0_control | _GEN_64; // @[LoopBlock.scala 903:56]
  assign _GEN_149 = loop_back_R_0_control | _GEN_66; // @[LoopBlock.scala 903:56]
  assign _GEN_150 = loop_back_R_0_control | _GEN_68; // @[LoopBlock.scala 903:56]
  assign _GEN_151 = loop_back_R_0_control | _GEN_70; // @[LoopBlock.scala 903:56]
  assign _GEN_152 = loop_back_R_0_control | _GEN_72; // @[LoopBlock.scala 903:56]
  assign _GEN_153 = loop_back_R_0_control | _GEN_74; // @[LoopBlock.scala 903:56]
  assign _T_101 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_4_ready = ~ in_live_in_valid_R_4; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_5_ready = ~ in_live_in_valid_R_5; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_6_ready = ~ in_live_in_valid_R_6; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_7_ready = ~ in_live_in_valid_R_7; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_8_ready = ~ in_live_in_valid_R_8; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field8_0_valid = out_live_in_valid_R_8_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field8_0_bits_taskID = in_live_in_R_8_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_bits_data = in_live_in_R_8_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_1_valid = out_live_in_valid_R_8_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field8_1_bits_data = in_live_in_R_8_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_valid = out_live_in_valid_R_7_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field7_0_bits_data = in_live_in_R_7_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_valid = out_live_in_valid_R_6_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field6_0_bits_data = in_live_in_R_6_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field5_0_bits_taskID = in_live_in_R_5_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_0_bits_taskID = in_live_in_R_4_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
  assign _GEN_454 = _T_60 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_455 = _GEN_454 & _T_73; // @[LoopBlock.scala 932:19]
  assign _GEN_456 = _GEN_455 & _T_85; // @[LoopBlock.scala 932:19]
  assign _GEN_457 = _GEN_456 & loop_back_R_0_control; // @[LoopBlock.scala 932:19]
  assign _GEN_461 = loop_back_R_0_control == 1'h0; // @[LoopBlock.scala 950:19]
  assign _GEN_462 = _GEN_456 & _GEN_461; // @[LoopBlock.scala 950:19]
  assign _GEN_463 = _GEN_462 & loop_finish_R_0_control; // @[LoopBlock.scala 950:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_4_taskID = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_4_data = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_R_5_taskID = _RAND_15[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_R_5_data = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_R_6_data = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_R_7_data = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_live_in_R_8_taskID = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_live_in_R_8_data = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  in_live_in_valid_R_6 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  in_live_in_valid_R_7 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  in_live_in_valid_R_8 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_30[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  out_live_in_valid_R_6_0 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  out_live_in_valid_R_7_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  out_live_in_valid_R_8_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  out_live_in_valid_R_8_1 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  out_live_in_fire_R_6_0 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  out_live_in_fire_R_7_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  out_live_in_fire_R_8_0 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  out_live_in_fire_R_8_1 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_54[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_57[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_60[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  state = _RAND_64[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_60) begin
        if (_T_21) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_73) begin
          if (_T_21) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_21) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_21) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_21) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_73) begin
          if (_T_21) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_21) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_21) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_60) begin
        enable_valid_R <= _GEN_3;
      end else begin
        if (_T_73) begin
          enable_valid_R <= _GEN_3;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_3;
            end
          end else begin
            enable_valid_R <= _GEN_3;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else begin
      if (_T_60) begin
        if (_T_23) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_23) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_23) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_23) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_23) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_23) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_23) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_23) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        loop_back_valid_R_0 <= _GEN_6;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_25) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_25) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_25) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_25) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_7;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        loop_finish_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_60) begin
        if (_T_27) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_73) begin
          if (_T_27) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_27) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_27) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_60) begin
        if (_T_29) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_73) begin
          if (_T_29) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_29) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_29) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_60) begin
        if (_T_31) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_73) begin
          if (_T_31) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_31) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_31) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_60) begin
        if (_T_33) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_73) begin
          if (_T_33) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_33) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_33) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_taskID <= 5'h0;
    end else begin
      if (_T_60) begin
        if (_T_35) begin
          in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
        end
      end else begin
        if (_T_73) begin
          if (_T_35) begin
            in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_taskID <= 5'h0;
            end else begin
              if (_T_35) begin
                in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
              end
            end
          end else begin
            if (_T_35) begin
              in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_data <= 32'h0;
    end else begin
      if (_T_60) begin
        if (_T_35) begin
          in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
        end
      end else begin
        if (_T_73) begin
          if (_T_35) begin
            in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_data <= 32'h0;
            end else begin
              if (_T_35) begin
                in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
              end
            end
          end else begin
            if (_T_35) begin
              in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_taskID <= 5'h0;
    end else begin
      if (_T_60) begin
        if (_T_37) begin
          in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
        end
      end else begin
        if (_T_73) begin
          if (_T_37) begin
            in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_taskID <= 5'h0;
            end else begin
              if (_T_37) begin
                in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
              end
            end
          end else begin
            if (_T_37) begin
              in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_data <= 32'h0;
    end else begin
      if (_T_60) begin
        if (_T_37) begin
          in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
        end
      end else begin
        if (_T_73) begin
          if (_T_37) begin
            in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_data <= 32'h0;
            end else begin
              if (_T_37) begin
                in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
              end
            end
          end else begin
            if (_T_37) begin
              in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_data <= 32'h0;
    end else begin
      if (_T_60) begin
        if (_T_39) begin
          in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
        end
      end else begin
        if (_T_73) begin
          if (_T_39) begin
            in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_data <= 32'h0;
            end else begin
              if (_T_39) begin
                in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
              end
            end
          end else begin
            if (_T_39) begin
              in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_data <= 32'h0;
    end else begin
      if (_T_60) begin
        if (_T_41) begin
          in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
        end
      end else begin
        if (_T_73) begin
          if (_T_41) begin
            in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_data <= 32'h0;
            end else begin
              if (_T_41) begin
                in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
              end
            end
          end else begin
            if (_T_41) begin
              in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_taskID <= 5'h0;
    end else begin
      if (_T_60) begin
        if (_T_43) begin
          in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
        end
      end else begin
        if (_T_73) begin
          if (_T_43) begin
            in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_taskID <= 5'h0;
            end else begin
              if (_T_43) begin
                in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
              end
            end
          end else begin
            if (_T_43) begin
              in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_data <= 32'h0;
    end else begin
      if (_T_60) begin
        if (_T_43) begin
          in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
        end
      end else begin
        if (_T_73) begin
          if (_T_43) begin
            in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_data <= 32'h0;
            end else begin
              if (_T_43) begin
                in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
              end
            end
          end else begin
            if (_T_43) begin
              in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_live_in_valid_R_0 <= _GEN_13;
      end else begin
        if (_T_73) begin
          in_live_in_valid_R_0 <= _GEN_13;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              in_live_in_valid_R_0 <= _GEN_13;
            end
          end else begin
            in_live_in_valid_R_0 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_live_in_valid_R_1 <= _GEN_17;
      end else begin
        if (_T_73) begin
          in_live_in_valid_R_1 <= _GEN_17;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              in_live_in_valid_R_1 <= _GEN_17;
            end
          end else begin
            in_live_in_valid_R_1 <= _GEN_17;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_live_in_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_73) begin
          in_live_in_valid_R_2 <= _GEN_21;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              in_live_in_valid_R_2 <= _GEN_21;
            end
          end else begin
            in_live_in_valid_R_2 <= _GEN_21;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_live_in_valid_R_3 <= _GEN_25;
      end else begin
        if (_T_73) begin
          in_live_in_valid_R_3 <= _GEN_25;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              in_live_in_valid_R_3 <= _GEN_25;
            end
          end else begin
            in_live_in_valid_R_3 <= _GEN_25;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_live_in_valid_R_4 <= _GEN_29;
      end else begin
        if (_T_73) begin
          in_live_in_valid_R_4 <= _GEN_29;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_4 <= 1'h0;
            end else begin
              in_live_in_valid_R_4 <= _GEN_29;
            end
          end else begin
            in_live_in_valid_R_4 <= _GEN_29;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_live_in_valid_R_5 <= _GEN_33;
      end else begin
        if (_T_73) begin
          in_live_in_valid_R_5 <= _GEN_33;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_5 <= 1'h0;
            end else begin
              in_live_in_valid_R_5 <= _GEN_33;
            end
          end else begin
            in_live_in_valid_R_5 <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_6 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_live_in_valid_R_6 <= _GEN_37;
      end else begin
        if (_T_73) begin
          in_live_in_valid_R_6 <= _GEN_37;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_6 <= 1'h0;
            end else begin
              in_live_in_valid_R_6 <= _GEN_37;
            end
          end else begin
            in_live_in_valid_R_6 <= _GEN_37;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_7 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_live_in_valid_R_7 <= _GEN_41;
      end else begin
        if (_T_73) begin
          in_live_in_valid_R_7 <= _GEN_41;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_7 <= 1'h0;
            end else begin
              in_live_in_valid_R_7 <= _GEN_41;
            end
          end else begin
            in_live_in_valid_R_7 <= _GEN_41;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_8 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_live_in_valid_R_8 <= _GEN_45;
      end else begin
        if (_T_73) begin
          in_live_in_valid_R_8 <= _GEN_45;
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_8 <= 1'h0;
            end else begin
              in_live_in_valid_R_8 <= _GEN_45;
            end
          end else begin
            in_live_in_valid_R_8 <= _GEN_45;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_45) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_45) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        in_carry_in_valid_R_0 <= _GEN_49;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_49;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_49;
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_49;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_49;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_0_0 <= _GEN_76;
        end else begin
          if (_T_49) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_0_0 <= _GEN_143;
          end else begin
            if (_T_49) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_49) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_1_0 <= _GEN_77;
        end else begin
          if (_T_50) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_1_0 <= _GEN_144;
          end else begin
            if (_T_50) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_50) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_2_0 <= _GEN_78;
        end else begin
          if (_T_51) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_2_0 <= _GEN_145;
          end else begin
            if (_T_51) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_51) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_3_0 <= _GEN_79;
        end else begin
          if (_T_52) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_3_0 <= _GEN_146;
          end else begin
            if (_T_52) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_52) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_4_0 <= _GEN_80;
        end else begin
          if (_T_53) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_4_0 <= _GEN_147;
          end else begin
            if (_T_53) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_53) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_5_0 <= _GEN_81;
        end else begin
          if (_T_54) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_5_0 <= _GEN_148;
          end else begin
            if (_T_54) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_54) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_6_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_6_0 <= _GEN_82;
        end else begin
          if (_T_55) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_6_0 <= _GEN_149;
          end else begin
            if (_T_55) begin
              out_live_in_valid_R_6_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_55) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_7_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_7_0 <= _GEN_83;
        end else begin
          if (_T_56) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_7_0 <= _GEN_150;
          end else begin
            if (_T_56) begin
              out_live_in_valid_R_7_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_56) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_8_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_8_0 <= _GEN_84;
        end else begin
          if (_T_57) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_8_0 <= _GEN_151;
          end else begin
            if (_T_57) begin
              out_live_in_valid_R_8_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_57) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_8_1 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_live_in_valid_R_8_1 <= _GEN_85;
        end else begin
          if (_T_58) begin
            out_live_in_valid_R_8_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_live_in_valid_R_8_1 <= _GEN_152;
          end else begin
            if (_T_58) begin
              out_live_in_valid_R_8_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_58) begin
            out_live_in_valid_R_8_1 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_0_0 <= _GEN_55;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_0 <= _GEN_55;
            end
          end else begin
            out_live_in_fire_R_0_0 <= _GEN_55;
          end
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_55;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_1_0 <= _GEN_57;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_0 <= _GEN_57;
            end
          end else begin
            out_live_in_fire_R_1_0 <= _GEN_57;
          end
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_57;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_2_0 <= _GEN_59;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_2_0 <= _GEN_59;
            end
          end else begin
            out_live_in_fire_R_2_0 <= _GEN_59;
          end
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_59;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_3_0 <= _GEN_61;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_3_0 <= _GEN_61;
            end
          end else begin
            out_live_in_fire_R_3_0 <= _GEN_61;
          end
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_61;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_4_0 <= _GEN_63;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_4_0 <= _GEN_63;
            end
          end else begin
            out_live_in_fire_R_4_0 <= _GEN_63;
          end
        end else begin
          out_live_in_fire_R_4_0 <= _GEN_63;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_5_0 <= _GEN_65;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_5_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_5_0 <= _GEN_65;
            end
          end else begin
            out_live_in_fire_R_5_0 <= _GEN_65;
          end
        end else begin
          out_live_in_fire_R_5_0 <= _GEN_65;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_6_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_6_0 <= _GEN_67;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_6_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_6_0 <= _GEN_67;
            end
          end else begin
            out_live_in_fire_R_6_0 <= _GEN_67;
          end
        end else begin
          out_live_in_fire_R_6_0 <= _GEN_67;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_7_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_7_0 <= _GEN_69;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_7_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_7_0 <= _GEN_69;
            end
          end else begin
            out_live_in_fire_R_7_0 <= _GEN_69;
          end
        end else begin
          out_live_in_fire_R_7_0 <= _GEN_69;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_8_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_8_0 <= _GEN_71;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_8_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_8_0 <= _GEN_71;
            end
          end else begin
            out_live_in_fire_R_8_0 <= _GEN_71;
          end
        end else begin
          out_live_in_fire_R_8_0 <= _GEN_71;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_8_1 <= 1'h0;
    end else begin
      if (_T_60) begin
        out_live_in_fire_R_8_1 <= _GEN_73;
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_8_1 <= 1'h0;
            end else begin
              out_live_in_fire_R_8_1 <= _GEN_73;
            end
          end else begin
            out_live_in_fire_R_8_1 <= _GEN_73;
          end
        end else begin
          out_live_in_fire_R_8_1 <= _GEN_73;
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          out_carry_out_valid_R_0_0 <= _GEN_86;
        end else begin
          if (_T_59) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            out_carry_out_valid_R_0_0 <= _GEN_153;
          end else begin
            if (_T_59) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_59) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          active_loop_start_R_control <= _GEN_87;
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          active_loop_start_valid_R <= _GEN_89;
        end else begin
          if (_T_46) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            active_loop_start_valid_R <= _GEN_128;
          end else begin
            if (_T_46) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_46) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            active_loop_back_R_control <= _GEN_129;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          active_loop_back_valid_R <= _GEN_92;
        end else begin
          if (_T_47) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            active_loop_back_valid_R <= _GEN_131;
          end else begin
            if (_T_47) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_47) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 5'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          loop_exit_R_0_control <= _GEN_94;
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (!(loop_back_R_0_control)) begin
              loop_exit_R_0_control <= _GEN_123;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          if (enable_R_control) begin
            if (_T_48) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_48) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              if (_T_48) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              loop_exit_valid_R_0 <= _GEN_118;
            end
          end else begin
            if (_T_48) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_52;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_53;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_60) begin
        if (_T_69) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_73) begin
          if (_T_85) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_101) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_457 & _T_93) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_3: Restarted fired @ %d\n",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 932:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_463 & _T_93) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_3: Output fired @ %d ",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 950:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_463 & _T_93) begin
          $fwrite(32'h80000002,"\n"); // @[LoopBlock.scala 955:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [4:0]  io_InLiveIn_3_bits_taskID,
  input  [31:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [4:0]  io_InLiveIn_4_bits_taskID,
  input  [31:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input  [31:0] io_InLiveIn_5_bits_data,
  output        io_InLiveIn_6_ready,
  input         io_InLiveIn_6_valid,
  input  [31:0] io_InLiveIn_6_bits_data,
  output        io_InLiveIn_7_ready,
  input         io_InLiveIn_7_valid,
  input  [4:0]  io_InLiveIn_7_bits_taskID,
  input  [31:0] io_InLiveIn_7_bits_data,
  output        io_InLiveIn_8_ready,
  input         io_InLiveIn_8_valid,
  input  [4:0]  io_InLiveIn_8_bits_taskID,
  input  [31:0] io_InLiveIn_8_bits_data,
  output        io_InLiveIn_9_ready,
  input         io_InLiveIn_9_valid,
  input  [31:0] io_InLiveIn_9_bits_data,
  output        io_InLiveIn_10_ready,
  input         io_InLiveIn_10_valid,
  input  [4:0]  io_InLiveIn_10_bits_taskID,
  input  [31:0] io_InLiveIn_10_bits_data,
  output        io_InLiveIn_11_ready,
  input         io_InLiveIn_11_valid,
  input  [31:0] io_InLiveIn_11_bits_data,
  input         io_OutLiveIn_field11_0_ready,
  output        io_OutLiveIn_field11_0_valid,
  output [31:0] io_OutLiveIn_field11_0_bits_data,
  input         io_OutLiveIn_field10_0_ready,
  output        io_OutLiveIn_field10_0_valid,
  output [4:0]  io_OutLiveIn_field10_0_bits_taskID,
  output [31:0] io_OutLiveIn_field10_0_bits_data,
  input         io_OutLiveIn_field10_1_ready,
  output        io_OutLiveIn_field10_1_valid,
  output [31:0] io_OutLiveIn_field10_1_bits_data,
  input         io_OutLiveIn_field9_0_ready,
  output        io_OutLiveIn_field9_0_valid,
  output [31:0] io_OutLiveIn_field9_0_bits_data,
  input         io_OutLiveIn_field8_0_ready,
  output        io_OutLiveIn_field8_0_valid,
  output [4:0]  io_OutLiveIn_field8_0_bits_taskID,
  output [31:0] io_OutLiveIn_field8_0_bits_data,
  input         io_OutLiveIn_field7_0_ready,
  output        io_OutLiveIn_field7_0_valid,
  output [4:0]  io_OutLiveIn_field7_0_bits_taskID,
  output [31:0] io_OutLiveIn_field7_0_bits_data,
  input         io_OutLiveIn_field6_0_ready,
  output        io_OutLiveIn_field6_0_valid,
  output [31:0] io_OutLiveIn_field6_0_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output [31:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [4:0]  io_OutLiveIn_field4_0_bits_taskID,
  output [31:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [4:0]  io_OutLiveIn_field3_0_bits_taskID,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_2;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_3;
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_5;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_6;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_7;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_8;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [4:0] in_live_in_R_3_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [4:0] in_live_in_R_4_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg [31:0] in_live_in_R_4_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_15;
  reg [31:0] in_live_in_R_5_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_16;
  reg [31:0] in_live_in_R_6_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_17;
  reg [4:0] in_live_in_R_7_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_18;
  reg [31:0] in_live_in_R_7_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_19;
  reg [4:0] in_live_in_R_8_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_20;
  reg [31:0] in_live_in_R_8_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_21;
  reg [31:0] in_live_in_R_9_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_22;
  reg [4:0] in_live_in_R_10_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_23;
  reg [31:0] in_live_in_R_10_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_24;
  reg [31:0] in_live_in_R_11_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_25;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_26;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_27;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_28;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_29;
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_30;
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_31;
  reg  in_live_in_valid_R_6; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_32;
  reg  in_live_in_valid_R_7; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_33;
  reg  in_live_in_valid_R_8; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_34;
  reg  in_live_in_valid_R_9; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_35;
  reg  in_live_in_valid_R_10; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_36;
  reg  in_live_in_valid_R_11; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_37;
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_38;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_39;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_40;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_41;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_42;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_43;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_44;
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_45;
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_46;
  reg  out_live_in_valid_R_6_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_47;
  reg  out_live_in_valid_R_7_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_48;
  reg  out_live_in_valid_R_8_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_49;
  reg  out_live_in_valid_R_9_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_50;
  reg  out_live_in_valid_R_10_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_51;
  reg  out_live_in_valid_R_10_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_52;
  reg  out_live_in_valid_R_11_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_53;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_54;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_55;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_56;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_57;
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_58;
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_59;
  reg  out_live_in_fire_R_6_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_60;
  reg  out_live_in_fire_R_7_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_61;
  reg  out_live_in_fire_R_8_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_62;
  reg  out_live_in_fire_R_9_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_63;
  reg  out_live_in_fire_R_10_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_64;
  reg  out_live_in_fire_R_10_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_65;
  reg  out_live_in_fire_R_11_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_66;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_67;
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_68;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_69;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_70;
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_71;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_72;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_73;
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_74;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_75;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_76;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_77;
  wire  _T_24; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_26; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[LoopBlock.scala 603:33]
  wire [4:0] _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_28; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_32; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_34; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_36; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_38; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[LoopBlock.scala 623:33]
  wire  _T_40; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[LoopBlock.scala 623:33]
  wire  _T_42; // @[Decoupled.scala 40:37]
  wire  _GEN_37; // @[LoopBlock.scala 623:33]
  wire  _T_44; // @[Decoupled.scala 40:37]
  wire  _GEN_41; // @[LoopBlock.scala 623:33]
  wire  _T_46; // @[Decoupled.scala 40:37]
  wire  _GEN_45; // @[LoopBlock.scala 623:33]
  wire  _T_48; // @[Decoupled.scala 40:37]
  wire  _GEN_49; // @[LoopBlock.scala 623:33]
  wire  _T_50; // @[Decoupled.scala 40:37]
  wire  _GEN_53; // @[LoopBlock.scala 623:33]
  wire  _T_52; // @[Decoupled.scala 40:37]
  wire  _GEN_57; // @[LoopBlock.scala 623:33]
  wire  _T_54; // @[Decoupled.scala 40:37]
  wire  _GEN_61; // @[LoopBlock.scala 641:37]
  wire  _T_55; // @[Decoupled.scala 40:37]
  wire  _GEN_62; // @[LoopBlock.scala 704:39]
  wire  _T_56; // @[Decoupled.scala 40:37]
  wire  _GEN_63; // @[LoopBlock.scala 708:38]
  wire  _T_57; // @[Decoupled.scala 40:37]
  wire  _GEN_64; // @[LoopBlock.scala 713:33]
  wire  _GEN_65; // @[LoopBlock.scala 713:33]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire  _GEN_66; // @[LoopBlock.scala 722:57]
  wire  _GEN_67; // @[LoopBlock.scala 722:57]
  wire  _T_59; // @[Decoupled.scala 40:37]
  wire  _GEN_68; // @[LoopBlock.scala 722:57]
  wire  _GEN_69; // @[LoopBlock.scala 722:57]
  wire  _T_60; // @[Decoupled.scala 40:37]
  wire  _GEN_70; // @[LoopBlock.scala 722:57]
  wire  _GEN_71; // @[LoopBlock.scala 722:57]
  wire  _T_61; // @[Decoupled.scala 40:37]
  wire  _GEN_72; // @[LoopBlock.scala 722:57]
  wire  _GEN_73; // @[LoopBlock.scala 722:57]
  wire  _T_62; // @[Decoupled.scala 40:37]
  wire  _GEN_74; // @[LoopBlock.scala 722:57]
  wire  _GEN_75; // @[LoopBlock.scala 722:57]
  wire  _T_63; // @[Decoupled.scala 40:37]
  wire  _GEN_76; // @[LoopBlock.scala 722:57]
  wire  _GEN_77; // @[LoopBlock.scala 722:57]
  wire  _T_64; // @[Decoupled.scala 40:37]
  wire  _GEN_78; // @[LoopBlock.scala 722:57]
  wire  _GEN_79; // @[LoopBlock.scala 722:57]
  wire  _T_65; // @[Decoupled.scala 40:37]
  wire  _GEN_80; // @[LoopBlock.scala 722:57]
  wire  _GEN_81; // @[LoopBlock.scala 722:57]
  wire  _T_66; // @[Decoupled.scala 40:37]
  wire  _GEN_82; // @[LoopBlock.scala 722:57]
  wire  _GEN_83; // @[LoopBlock.scala 722:57]
  wire  _T_67; // @[Decoupled.scala 40:37]
  wire  _GEN_84; // @[LoopBlock.scala 722:57]
  wire  _GEN_85; // @[LoopBlock.scala 722:57]
  wire  _T_68; // @[Decoupled.scala 40:37]
  wire  _GEN_86; // @[LoopBlock.scala 722:57]
  wire  _GEN_87; // @[LoopBlock.scala 722:57]
  wire  _T_69; // @[Decoupled.scala 40:37]
  wire  _GEN_88; // @[LoopBlock.scala 722:57]
  wire  _GEN_89; // @[LoopBlock.scala 722:57]
  wire  _T_70; // @[Decoupled.scala 40:37]
  wire  _GEN_90; // @[LoopBlock.scala 722:57]
  wire  _GEN_91; // @[LoopBlock.scala 722:57]
  wire  _T_71; // @[Decoupled.scala 40:37]
  wire  _GEN_92; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_78;
  wire  _T_72; // @[Conditional.scala 37:30]
  wire  _T_73; // @[LoopBlock.scala 765:35]
  wire  _T_74; // @[LoopBlock.scala 765:35]
  wire  _T_75; // @[LoopBlock.scala 765:35]
  wire  _T_76; // @[LoopBlock.scala 765:35]
  wire  _T_77; // @[LoopBlock.scala 765:35]
  wire  _T_78; // @[LoopBlock.scala 765:35]
  wire  _T_79; // @[LoopBlock.scala 765:35]
  wire  _T_80; // @[LoopBlock.scala 765:35]
  wire  _T_81; // @[LoopBlock.scala 765:35]
  wire  _T_82; // @[LoopBlock.scala 765:35]
  wire  _T_83; // @[LoopBlock.scala 765:35]
  wire  _T_84; // @[LoopBlock.scala 869:28]
  wire  _GEN_94; // @[LoopBlock.scala 870:26]
  wire  _GEN_95; // @[LoopBlock.scala 870:26]
  wire  _GEN_96; // @[LoopBlock.scala 870:26]
  wire  _GEN_97; // @[LoopBlock.scala 870:26]
  wire  _GEN_98; // @[LoopBlock.scala 870:26]
  wire  _GEN_99; // @[LoopBlock.scala 870:26]
  wire  _GEN_100; // @[LoopBlock.scala 870:26]
  wire  _GEN_101; // @[LoopBlock.scala 870:26]
  wire  _GEN_102; // @[LoopBlock.scala 870:26]
  wire  _GEN_103; // @[LoopBlock.scala 870:26]
  wire  _GEN_104; // @[LoopBlock.scala 870:26]
  wire  _GEN_105; // @[LoopBlock.scala 870:26]
  wire  _GEN_106; // @[LoopBlock.scala 870:26]
  wire  _GEN_107; // @[LoopBlock.scala 870:26]
  wire  _GEN_108; // @[LoopBlock.scala 870:26]
  wire  _GEN_110; // @[LoopBlock.scala 870:26]
  wire  _GEN_113; // @[LoopBlock.scala 870:26]
  wire  _GEN_115; // @[LoopBlock.scala 870:26]
  wire  _T_88; // @[Conditional.scala 37:30]
  wire  _T_89; // @[LoopBlock.scala 898:30]
  wire  _T_91; // @[LoopBlock.scala 825:65]
  wire  _T_92; // @[LoopBlock.scala 828:26]
  wire  _T_93; // @[LoopBlock.scala 828:26]
  wire  _T_94; // @[LoopBlock.scala 828:26]
  wire  _T_95; // @[LoopBlock.scala 828:26]
  wire  _T_96; // @[LoopBlock.scala 828:26]
  wire  _T_97; // @[LoopBlock.scala 828:26]
  wire  _T_98; // @[LoopBlock.scala 828:26]
  wire  _T_99; // @[LoopBlock.scala 828:26]
  wire  _T_100; // @[LoopBlock.scala 828:26]
  wire  _T_101; // @[LoopBlock.scala 828:26]
  wire  _T_102; // @[LoopBlock.scala 828:26]
  wire  _T_103; // @[LoopBlock.scala 899:29]
  wire  _T_110; // @[LoopBlock.scala 932:19]
  wire  _T_111; // @[LoopBlock.scala 932:19]
  wire  _GEN_142; // @[LoopBlock.scala 936:64]
  wire  _GEN_145; // @[LoopBlock.scala 936:64]
  wire  _GEN_147; // @[LoopBlock.scala 936:64]
  wire  _GEN_152; // @[LoopBlock.scala 903:56]
  wire  _GEN_153; // @[LoopBlock.scala 903:56]
  wire  _GEN_155; // @[LoopBlock.scala 903:56]
  wire  _GEN_170; // @[LoopBlock.scala 903:56]
  wire  _GEN_171; // @[LoopBlock.scala 903:56]
  wire  _GEN_172; // @[LoopBlock.scala 903:56]
  wire  _GEN_173; // @[LoopBlock.scala 903:56]
  wire  _GEN_174; // @[LoopBlock.scala 903:56]
  wire  _GEN_175; // @[LoopBlock.scala 903:56]
  wire  _GEN_176; // @[LoopBlock.scala 903:56]
  wire  _GEN_177; // @[LoopBlock.scala 903:56]
  wire  _GEN_178; // @[LoopBlock.scala 903:56]
  wire  _GEN_179; // @[LoopBlock.scala 903:56]
  wire  _GEN_180; // @[LoopBlock.scala 903:56]
  wire  _GEN_181; // @[LoopBlock.scala 903:56]
  wire  _GEN_182; // @[LoopBlock.scala 903:56]
  wire  _GEN_183; // @[LoopBlock.scala 903:56]
  wire  _T_119; // @[Conditional.scala 37:30]
  wire  _GEN_550; // @[LoopBlock.scala 932:19]
  wire  _GEN_551; // @[LoopBlock.scala 932:19]
  wire  _GEN_552; // @[LoopBlock.scala 932:19]
  wire  _GEN_553; // @[LoopBlock.scala 932:19]
  wire  _GEN_557; // @[LoopBlock.scala 950:19]
  wire  _GEN_558; // @[LoopBlock.scala 950:19]
  wire  _GEN_559; // @[LoopBlock.scala 950:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_24 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_24 | enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_26 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_26 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_26 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_26 | loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_28 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_28 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_28 | loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_30 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_30 | in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_32 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_32 | in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_34 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_34 | in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_36 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_36 | in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_38 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_38 | in_live_in_valid_R_4; // @[LoopBlock.scala 623:33]
  assign _T_40 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_40 | in_live_in_valid_R_5; // @[LoopBlock.scala 623:33]
  assign _T_42 = io_InLiveIn_6_ready & io_InLiveIn_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_37 = _T_42 | in_live_in_valid_R_6; // @[LoopBlock.scala 623:33]
  assign _T_44 = io_InLiveIn_7_ready & io_InLiveIn_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_41 = _T_44 | in_live_in_valid_R_7; // @[LoopBlock.scala 623:33]
  assign _T_46 = io_InLiveIn_8_ready & io_InLiveIn_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_45 = _T_46 | in_live_in_valid_R_8; // @[LoopBlock.scala 623:33]
  assign _T_48 = io_InLiveIn_9_ready & io_InLiveIn_9_valid; // @[Decoupled.scala 40:37]
  assign _GEN_49 = _T_48 | in_live_in_valid_R_9; // @[LoopBlock.scala 623:33]
  assign _T_50 = io_InLiveIn_10_ready & io_InLiveIn_10_valid; // @[Decoupled.scala 40:37]
  assign _GEN_53 = _T_50 | in_live_in_valid_R_10; // @[LoopBlock.scala 623:33]
  assign _T_52 = io_InLiveIn_11_ready & io_InLiveIn_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_57 = _T_52 | in_live_in_valid_R_11; // @[LoopBlock.scala 623:33]
  assign _T_54 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_61 = _T_54 | in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_55 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  assign _GEN_62 = _T_55 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_56 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  assign _GEN_63 = _T_56 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_57 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_64 = _T_57 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_65 = _T_57 | loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_58 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_66 = _T_58 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_67 = _T_58 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_59 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_68 = _T_59 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_69 = _T_59 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_60 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_70 = _T_60 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_71 = _T_60 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_61 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_72 = _T_61 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_73 = _T_61 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_62 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_74 = _T_62 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 722:57]
  assign _GEN_75 = _T_62 | out_live_in_fire_R_4_0; // @[LoopBlock.scala 722:57]
  assign _T_63 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_76 = _T_63 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 722:57]
  assign _GEN_77 = _T_63 | out_live_in_fire_R_5_0; // @[LoopBlock.scala 722:57]
  assign _T_64 = io_OutLiveIn_field6_0_ready & io_OutLiveIn_field6_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_78 = _T_64 ? 1'h0 : out_live_in_valid_R_6_0; // @[LoopBlock.scala 722:57]
  assign _GEN_79 = _T_64 | out_live_in_fire_R_6_0; // @[LoopBlock.scala 722:57]
  assign _T_65 = io_OutLiveIn_field7_0_ready & io_OutLiveIn_field7_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_80 = _T_65 ? 1'h0 : out_live_in_valid_R_7_0; // @[LoopBlock.scala 722:57]
  assign _GEN_81 = _T_65 | out_live_in_fire_R_7_0; // @[LoopBlock.scala 722:57]
  assign _T_66 = io_OutLiveIn_field8_0_ready & io_OutLiveIn_field8_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_82 = _T_66 ? 1'h0 : out_live_in_valid_R_8_0; // @[LoopBlock.scala 722:57]
  assign _GEN_83 = _T_66 | out_live_in_fire_R_8_0; // @[LoopBlock.scala 722:57]
  assign _T_67 = io_OutLiveIn_field9_0_ready & io_OutLiveIn_field9_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_84 = _T_67 ? 1'h0 : out_live_in_valid_R_9_0; // @[LoopBlock.scala 722:57]
  assign _GEN_85 = _T_67 | out_live_in_fire_R_9_0; // @[LoopBlock.scala 722:57]
  assign _T_68 = io_OutLiveIn_field10_0_ready & io_OutLiveIn_field10_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_86 = _T_68 ? 1'h0 : out_live_in_valid_R_10_0; // @[LoopBlock.scala 722:57]
  assign _GEN_87 = _T_68 | out_live_in_fire_R_10_0; // @[LoopBlock.scala 722:57]
  assign _T_69 = io_OutLiveIn_field10_1_ready & io_OutLiveIn_field10_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_88 = _T_69 ? 1'h0 : out_live_in_valid_R_10_1; // @[LoopBlock.scala 722:57]
  assign _GEN_89 = _T_69 | out_live_in_fire_R_10_1; // @[LoopBlock.scala 722:57]
  assign _T_70 = io_OutLiveIn_field11_0_ready & io_OutLiveIn_field11_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_90 = _T_70 ? 1'h0 : out_live_in_valid_R_11_0; // @[LoopBlock.scala 722:57]
  assign _GEN_91 = _T_70 | out_live_in_fire_R_11_0; // @[LoopBlock.scala 722:57]
  assign _T_71 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_92 = _T_71 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_72 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_73 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_74 = _T_73 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_75 = _T_74 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_76 = _T_75 & in_live_in_valid_R_4; // @[LoopBlock.scala 765:35]
  assign _T_77 = _T_76 & in_live_in_valid_R_5; // @[LoopBlock.scala 765:35]
  assign _T_78 = _T_77 & in_live_in_valid_R_6; // @[LoopBlock.scala 765:35]
  assign _T_79 = _T_78 & in_live_in_valid_R_7; // @[LoopBlock.scala 765:35]
  assign _T_80 = _T_79 & in_live_in_valid_R_8; // @[LoopBlock.scala 765:35]
  assign _T_81 = _T_80 & in_live_in_valid_R_9; // @[LoopBlock.scala 765:35]
  assign _T_82 = _T_81 & in_live_in_valid_R_10; // @[LoopBlock.scala 765:35]
  assign _T_83 = _T_82 & in_live_in_valid_R_11; // @[LoopBlock.scala 765:35]
  assign _T_84 = _T_83 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_94 = enable_R_control | _GEN_66; // @[LoopBlock.scala 870:26]
  assign _GEN_95 = enable_R_control | _GEN_68; // @[LoopBlock.scala 870:26]
  assign _GEN_96 = enable_R_control | _GEN_70; // @[LoopBlock.scala 870:26]
  assign _GEN_97 = enable_R_control | _GEN_72; // @[LoopBlock.scala 870:26]
  assign _GEN_98 = enable_R_control | _GEN_74; // @[LoopBlock.scala 870:26]
  assign _GEN_99 = enable_R_control | _GEN_76; // @[LoopBlock.scala 870:26]
  assign _GEN_100 = enable_R_control | _GEN_78; // @[LoopBlock.scala 870:26]
  assign _GEN_101 = enable_R_control | _GEN_80; // @[LoopBlock.scala 870:26]
  assign _GEN_102 = enable_R_control | _GEN_82; // @[LoopBlock.scala 870:26]
  assign _GEN_103 = enable_R_control | _GEN_84; // @[LoopBlock.scala 870:26]
  assign _GEN_104 = enable_R_control | _GEN_86; // @[LoopBlock.scala 870:26]
  assign _GEN_105 = enable_R_control | _GEN_88; // @[LoopBlock.scala 870:26]
  assign _GEN_106 = enable_R_control | _GEN_90; // @[LoopBlock.scala 870:26]
  assign _GEN_107 = enable_R_control | _GEN_92; // @[LoopBlock.scala 870:26]
  assign _GEN_108 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_110 = enable_R_control | _GEN_62; // @[LoopBlock.scala 870:26]
  assign _GEN_113 = enable_R_control | _GEN_63; // @[LoopBlock.scala 870:26]
  assign _GEN_115 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 870:26]
  assign _T_88 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_89 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_91 = out_live_in_fire_R_10_0 & out_live_in_fire_R_10_1; // @[LoopBlock.scala 825:65]
  assign _T_92 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_93 = _T_92 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_94 = _T_93 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_95 = _T_94 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 828:26]
  assign _T_96 = _T_95 & out_live_in_fire_R_5_0; // @[LoopBlock.scala 828:26]
  assign _T_97 = _T_96 & out_live_in_fire_R_6_0; // @[LoopBlock.scala 828:26]
  assign _T_98 = _T_97 & out_live_in_fire_R_7_0; // @[LoopBlock.scala 828:26]
  assign _T_99 = _T_98 & out_live_in_fire_R_8_0; // @[LoopBlock.scala 828:26]
  assign _T_100 = _T_99 & out_live_in_fire_R_9_0; // @[LoopBlock.scala 828:26]
  assign _T_101 = _T_100 & _T_91; // @[LoopBlock.scala 828:26]
  assign _T_102 = _T_101 & out_live_in_fire_R_11_0; // @[LoopBlock.scala 828:26]
  assign _T_103 = _T_89 & _T_102; // @[LoopBlock.scala 899:29]
  assign _T_110 = $unsigned(reset); // @[LoopBlock.scala 932:19]
  assign _T_111 = _T_110 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_142 = loop_finish_R_0_control | _GEN_64; // @[LoopBlock.scala 936:64]
  assign _GEN_145 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_147 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_152 = loop_back_R_0_control | _GEN_62; // @[LoopBlock.scala 903:56]
  assign _GEN_153 = loop_back_R_0_control | _GEN_145; // @[LoopBlock.scala 903:56]
  assign _GEN_155 = loop_back_R_0_control | _GEN_63; // @[LoopBlock.scala 903:56]
  assign _GEN_170 = loop_back_R_0_control | _GEN_66; // @[LoopBlock.scala 903:56]
  assign _GEN_171 = loop_back_R_0_control | _GEN_68; // @[LoopBlock.scala 903:56]
  assign _GEN_172 = loop_back_R_0_control | _GEN_70; // @[LoopBlock.scala 903:56]
  assign _GEN_173 = loop_back_R_0_control | _GEN_72; // @[LoopBlock.scala 903:56]
  assign _GEN_174 = loop_back_R_0_control | _GEN_74; // @[LoopBlock.scala 903:56]
  assign _GEN_175 = loop_back_R_0_control | _GEN_76; // @[LoopBlock.scala 903:56]
  assign _GEN_176 = loop_back_R_0_control | _GEN_78; // @[LoopBlock.scala 903:56]
  assign _GEN_177 = loop_back_R_0_control | _GEN_80; // @[LoopBlock.scala 903:56]
  assign _GEN_178 = loop_back_R_0_control | _GEN_82; // @[LoopBlock.scala 903:56]
  assign _GEN_179 = loop_back_R_0_control | _GEN_84; // @[LoopBlock.scala 903:56]
  assign _GEN_180 = loop_back_R_0_control | _GEN_86; // @[LoopBlock.scala 903:56]
  assign _GEN_181 = loop_back_R_0_control | _GEN_88; // @[LoopBlock.scala 903:56]
  assign _GEN_182 = loop_back_R_0_control | _GEN_90; // @[LoopBlock.scala 903:56]
  assign _GEN_183 = loop_back_R_0_control | _GEN_92; // @[LoopBlock.scala 903:56]
  assign _T_119 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_4_ready = ~ in_live_in_valid_R_4; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_5_ready = ~ in_live_in_valid_R_5; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_6_ready = ~ in_live_in_valid_R_6; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_7_ready = ~ in_live_in_valid_R_7; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_8_ready = ~ in_live_in_valid_R_8; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_9_ready = ~ in_live_in_valid_R_9; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_10_ready = ~ in_live_in_valid_R_10; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_11_ready = ~ in_live_in_valid_R_11; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field11_0_valid = out_live_in_valid_R_11_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field11_0_bits_data = in_live_in_R_11_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_0_valid = out_live_in_valid_R_10_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_0_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_0_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_1_valid = out_live_in_valid_R_10_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_1_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field9_0_valid = out_live_in_valid_R_9_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field9_0_bits_data = in_live_in_R_9_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_valid = out_live_in_valid_R_8_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field8_0_bits_taskID = in_live_in_R_8_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_bits_data = in_live_in_R_8_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_valid = out_live_in_valid_R_7_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field7_0_bits_taskID = in_live_in_R_7_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_bits_data = in_live_in_R_7_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_valid = out_live_in_valid_R_6_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field6_0_bits_data = in_live_in_R_6_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_0_bits_taskID = in_live_in_R_4_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_taskID = in_live_in_R_3_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
  assign _GEN_550 = _T_72 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_551 = _GEN_550 & _T_88; // @[LoopBlock.scala 932:19]
  assign _GEN_552 = _GEN_551 & _T_103; // @[LoopBlock.scala 932:19]
  assign _GEN_553 = _GEN_552 & loop_back_R_0_control; // @[LoopBlock.scala 932:19]
  assign _GEN_557 = loop_back_R_0_control == 1'h0; // @[LoopBlock.scala 950:19]
  assign _GEN_558 = _GEN_552 & _GEN_557; // @[LoopBlock.scala 950:19]
  assign _GEN_559 = _GEN_558 & loop_finish_R_0_control; // @[LoopBlock.scala 950:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_3_taskID = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_4_taskID = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_R_4_data = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_R_5_data = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_R_6_data = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_R_7_taskID = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_live_in_R_7_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_live_in_R_8_taskID = _RAND_20[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_live_in_R_8_data = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_live_in_R_9_data = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_live_in_R_10_taskID = _RAND_23[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_live_in_R_10_data = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_live_in_R_11_data = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  in_live_in_valid_R_6 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  in_live_in_valid_R_7 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  in_live_in_valid_R_8 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  in_live_in_valid_R_9 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  in_live_in_valid_R_10 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  in_live_in_valid_R_11 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_38[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  out_live_in_valid_R_6_0 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  out_live_in_valid_R_7_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  out_live_in_valid_R_8_0 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  out_live_in_valid_R_9_0 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  out_live_in_valid_R_10_0 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  out_live_in_valid_R_10_1 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  out_live_in_valid_R_11_0 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  out_live_in_fire_R_6_0 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  out_live_in_fire_R_7_0 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  out_live_in_fire_R_8_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  out_live_in_fire_R_9_0 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  out_live_in_fire_R_10_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  out_live_in_fire_R_10_1 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  out_live_in_fire_R_11_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_68[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_71[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_74[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  state = _RAND_78[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_24) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_88) begin
          if (_T_24) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_24) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_24) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_24) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_88) begin
          if (_T_24) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_24) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_24) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_72) begin
        enable_valid_R <= _GEN_3;
      end else begin
        if (_T_88) begin
          enable_valid_R <= _GEN_3;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_3;
            end
          end else begin
            enable_valid_R <= _GEN_3;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_26) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_26) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_26) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_26) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_26) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_26) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_26) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_26) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        loop_back_valid_R_0 <= _GEN_6;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_28) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_28) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_28) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_28) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_7;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        loop_finish_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_30) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_30) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_30) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_30) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_32) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_32) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_32) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_32) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_34) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_34) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_34) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_34) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_36) begin
          in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
        end
      end else begin
        if (_T_88) begin
          if (_T_36) begin
            in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_taskID <= 5'h0;
            end else begin
              if (_T_36) begin
                in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
              end
            end
          end else begin
            if (_T_36) begin
              in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_36) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_36) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_36) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_36) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_38) begin
          in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
        end
      end else begin
        if (_T_88) begin
          if (_T_38) begin
            in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_taskID <= 5'h0;
            end else begin
              if (_T_38) begin
                in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
              end
            end
          end else begin
            if (_T_38) begin
              in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_38) begin
          in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_38) begin
            in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_data <= 32'h0;
            end else begin
              if (_T_38) begin
                in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
              end
            end
          end else begin
            if (_T_38) begin
              in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_40) begin
          in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_40) begin
            in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_data <= 32'h0;
            end else begin
              if (_T_40) begin
                in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
              end
            end
          end else begin
            if (_T_40) begin
              in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_42) begin
          in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_42) begin
            in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_data <= 32'h0;
            end else begin
              if (_T_42) begin
                in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
              end
            end
          end else begin
            if (_T_42) begin
              in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_44) begin
          in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
        end
      end else begin
        if (_T_88) begin
          if (_T_44) begin
            in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_taskID <= 5'h0;
            end else begin
              if (_T_44) begin
                in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
              end
            end
          end else begin
            if (_T_44) begin
              in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_44) begin
          in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_44) begin
            in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_data <= 32'h0;
            end else begin
              if (_T_44) begin
                in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
              end
            end
          end else begin
            if (_T_44) begin
              in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_46) begin
          in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
        end
      end else begin
        if (_T_88) begin
          if (_T_46) begin
            in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_taskID <= 5'h0;
            end else begin
              if (_T_46) begin
                in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
              end
            end
          end else begin
            if (_T_46) begin
              in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_46) begin
          in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_46) begin
            in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_data <= 32'h0;
            end else begin
              if (_T_46) begin
                in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
              end
            end
          end else begin
            if (_T_46) begin
              in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_9_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_48) begin
          in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_48) begin
            in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_9_data <= 32'h0;
            end else begin
              if (_T_48) begin
                in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
              end
            end
          end else begin
            if (_T_48) begin
              in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_10_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_50) begin
          in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
        end
      end else begin
        if (_T_88) begin
          if (_T_50) begin
            in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_10_taskID <= 5'h0;
            end else begin
              if (_T_50) begin
                in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
              end
            end
          end else begin
            if (_T_50) begin
              in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_10_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_50) begin
          in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_50) begin
            in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_10_data <= 32'h0;
            end else begin
              if (_T_50) begin
                in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
              end
            end
          end else begin
            if (_T_50) begin
              in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_11_data <= 32'h0;
    end else begin
      if (_T_72) begin
        if (_T_52) begin
          in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
        end
      end else begin
        if (_T_88) begin
          if (_T_52) begin
            in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_11_data <= 32'h0;
            end else begin
              if (_T_52) begin
                in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
              end
            end
          end else begin
            if (_T_52) begin
              in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_0 <= _GEN_13;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_0 <= _GEN_13;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              in_live_in_valid_R_0 <= _GEN_13;
            end
          end else begin
            in_live_in_valid_R_0 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_1 <= _GEN_17;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_1 <= _GEN_17;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              in_live_in_valid_R_1 <= _GEN_17;
            end
          end else begin
            in_live_in_valid_R_1 <= _GEN_17;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_2 <= _GEN_21;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              in_live_in_valid_R_2 <= _GEN_21;
            end
          end else begin
            in_live_in_valid_R_2 <= _GEN_21;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_3 <= _GEN_25;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_3 <= _GEN_25;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              in_live_in_valid_R_3 <= _GEN_25;
            end
          end else begin
            in_live_in_valid_R_3 <= _GEN_25;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_4 <= _GEN_29;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_4 <= _GEN_29;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_4 <= 1'h0;
            end else begin
              in_live_in_valid_R_4 <= _GEN_29;
            end
          end else begin
            in_live_in_valid_R_4 <= _GEN_29;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_5 <= _GEN_33;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_5 <= _GEN_33;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_5 <= 1'h0;
            end else begin
              in_live_in_valid_R_5 <= _GEN_33;
            end
          end else begin
            in_live_in_valid_R_5 <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_6 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_6 <= _GEN_37;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_6 <= _GEN_37;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_6 <= 1'h0;
            end else begin
              in_live_in_valid_R_6 <= _GEN_37;
            end
          end else begin
            in_live_in_valid_R_6 <= _GEN_37;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_7 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_7 <= _GEN_41;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_7 <= _GEN_41;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_7 <= 1'h0;
            end else begin
              in_live_in_valid_R_7 <= _GEN_41;
            end
          end else begin
            in_live_in_valid_R_7 <= _GEN_41;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_8 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_8 <= _GEN_45;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_8 <= _GEN_45;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_8 <= 1'h0;
            end else begin
              in_live_in_valid_R_8 <= _GEN_45;
            end
          end else begin
            in_live_in_valid_R_8 <= _GEN_45;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_9 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_9 <= _GEN_49;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_9 <= _GEN_49;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_9 <= 1'h0;
            end else begin
              in_live_in_valid_R_9 <= _GEN_49;
            end
          end else begin
            in_live_in_valid_R_9 <= _GEN_49;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_10 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_10 <= _GEN_53;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_10 <= _GEN_53;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_10 <= 1'h0;
            end else begin
              in_live_in_valid_R_10 <= _GEN_53;
            end
          end else begin
            in_live_in_valid_R_10 <= _GEN_53;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_11 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_live_in_valid_R_11 <= _GEN_57;
      end else begin
        if (_T_88) begin
          in_live_in_valid_R_11 <= _GEN_57;
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_11 <= 1'h0;
            end else begin
              in_live_in_valid_R_11 <= _GEN_57;
            end
          end else begin
            in_live_in_valid_R_11 <= _GEN_57;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_54) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_54) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        in_carry_in_valid_R_0 <= _GEN_61;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_61;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_61;
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_61;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_61;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_0_0 <= _GEN_94;
        end else begin
          if (_T_58) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_0_0 <= _GEN_170;
          end else begin
            if (_T_58) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_58) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_1_0 <= _GEN_95;
        end else begin
          if (_T_59) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_1_0 <= _GEN_171;
          end else begin
            if (_T_59) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_59) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_2_0 <= _GEN_96;
        end else begin
          if (_T_60) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_2_0 <= _GEN_172;
          end else begin
            if (_T_60) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_60) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_3_0 <= _GEN_97;
        end else begin
          if (_T_61) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_3_0 <= _GEN_173;
          end else begin
            if (_T_61) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_61) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_4_0 <= _GEN_98;
        end else begin
          if (_T_62) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_4_0 <= _GEN_174;
          end else begin
            if (_T_62) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_62) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_5_0 <= _GEN_99;
        end else begin
          if (_T_63) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_5_0 <= _GEN_175;
          end else begin
            if (_T_63) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_63) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_6_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_6_0 <= _GEN_100;
        end else begin
          if (_T_64) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_6_0 <= _GEN_176;
          end else begin
            if (_T_64) begin
              out_live_in_valid_R_6_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_64) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_7_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_7_0 <= _GEN_101;
        end else begin
          if (_T_65) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_7_0 <= _GEN_177;
          end else begin
            if (_T_65) begin
              out_live_in_valid_R_7_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_65) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_8_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_8_0 <= _GEN_102;
        end else begin
          if (_T_66) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_8_0 <= _GEN_178;
          end else begin
            if (_T_66) begin
              out_live_in_valid_R_8_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_66) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_9_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_9_0 <= _GEN_103;
        end else begin
          if (_T_67) begin
            out_live_in_valid_R_9_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_9_0 <= _GEN_179;
          end else begin
            if (_T_67) begin
              out_live_in_valid_R_9_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_67) begin
            out_live_in_valid_R_9_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_10_0 <= _GEN_104;
        end else begin
          if (_T_68) begin
            out_live_in_valid_R_10_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_10_0 <= _GEN_180;
          end else begin
            if (_T_68) begin
              out_live_in_valid_R_10_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_68) begin
            out_live_in_valid_R_10_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_1 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_10_1 <= _GEN_105;
        end else begin
          if (_T_69) begin
            out_live_in_valid_R_10_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_10_1 <= _GEN_181;
          end else begin
            if (_T_69) begin
              out_live_in_valid_R_10_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_69) begin
            out_live_in_valid_R_10_1 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_11_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_live_in_valid_R_11_0 <= _GEN_106;
        end else begin
          if (_T_70) begin
            out_live_in_valid_R_11_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_live_in_valid_R_11_0 <= _GEN_182;
          end else begin
            if (_T_70) begin
              out_live_in_valid_R_11_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_70) begin
            out_live_in_valid_R_11_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_0_0 <= _GEN_67;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_0 <= _GEN_67;
            end
          end else begin
            out_live_in_fire_R_0_0 <= _GEN_67;
          end
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_67;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_1_0 <= _GEN_69;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_0 <= _GEN_69;
            end
          end else begin
            out_live_in_fire_R_1_0 <= _GEN_69;
          end
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_69;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_2_0 <= _GEN_71;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_2_0 <= _GEN_71;
            end
          end else begin
            out_live_in_fire_R_2_0 <= _GEN_71;
          end
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_71;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_3_0 <= _GEN_73;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_3_0 <= _GEN_73;
            end
          end else begin
            out_live_in_fire_R_3_0 <= _GEN_73;
          end
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_73;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_4_0 <= _GEN_75;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_4_0 <= _GEN_75;
            end
          end else begin
            out_live_in_fire_R_4_0 <= _GEN_75;
          end
        end else begin
          out_live_in_fire_R_4_0 <= _GEN_75;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_5_0 <= _GEN_77;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_5_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_5_0 <= _GEN_77;
            end
          end else begin
            out_live_in_fire_R_5_0 <= _GEN_77;
          end
        end else begin
          out_live_in_fire_R_5_0 <= _GEN_77;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_6_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_6_0 <= _GEN_79;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_6_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_6_0 <= _GEN_79;
            end
          end else begin
            out_live_in_fire_R_6_0 <= _GEN_79;
          end
        end else begin
          out_live_in_fire_R_6_0 <= _GEN_79;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_7_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_7_0 <= _GEN_81;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_7_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_7_0 <= _GEN_81;
            end
          end else begin
            out_live_in_fire_R_7_0 <= _GEN_81;
          end
        end else begin
          out_live_in_fire_R_7_0 <= _GEN_81;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_8_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_8_0 <= _GEN_83;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_8_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_8_0 <= _GEN_83;
            end
          end else begin
            out_live_in_fire_R_8_0 <= _GEN_83;
          end
        end else begin
          out_live_in_fire_R_8_0 <= _GEN_83;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_9_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_9_0 <= _GEN_85;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_9_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_9_0 <= _GEN_85;
            end
          end else begin
            out_live_in_fire_R_9_0 <= _GEN_85;
          end
        end else begin
          out_live_in_fire_R_9_0 <= _GEN_85;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_10_0 <= _GEN_87;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_0 <= _GEN_87;
            end
          end else begin
            out_live_in_fire_R_10_0 <= _GEN_87;
          end
        end else begin
          out_live_in_fire_R_10_0 <= _GEN_87;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_1 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_10_1 <= _GEN_89;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_1 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_1 <= _GEN_89;
            end
          end else begin
            out_live_in_fire_R_10_1 <= _GEN_89;
          end
        end else begin
          out_live_in_fire_R_10_1 <= _GEN_89;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_11_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        out_live_in_fire_R_11_0 <= _GEN_91;
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_11_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_11_0 <= _GEN_91;
            end
          end else begin
            out_live_in_fire_R_11_0 <= _GEN_91;
          end
        end else begin
          out_live_in_fire_R_11_0 <= _GEN_91;
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          out_carry_out_valid_R_0_0 <= _GEN_107;
        end else begin
          if (_T_71) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            out_carry_out_valid_R_0_0 <= _GEN_183;
          end else begin
            if (_T_71) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_71) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          active_loop_start_R_control <= _GEN_108;
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          active_loop_start_valid_R <= _GEN_110;
        end else begin
          if (_T_55) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            active_loop_start_valid_R <= _GEN_152;
          end else begin
            if (_T_55) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_55) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            active_loop_back_R_control <= _GEN_153;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          active_loop_back_valid_R <= _GEN_113;
        end else begin
          if (_T_56) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            active_loop_back_valid_R <= _GEN_155;
          end else begin
            if (_T_56) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_56) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 5'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          loop_exit_R_0_control <= _GEN_115;
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (!(loop_back_R_0_control)) begin
              loop_exit_R_0_control <= _GEN_147;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          if (enable_R_control) begin
            if (_T_57) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_57) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              if (_T_57) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              loop_exit_valid_R_0 <= _GEN_142;
            end
          end else begin
            if (_T_57) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_64;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_65;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_72) begin
        if (_T_84) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_88) begin
          if (_T_103) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_119) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_553 & _T_111) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_4: Restarted fired @ %d\n",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 932:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_559 & _T_111) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_4: Output fired @ %d ",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 950:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_559 & _T_111) begin
          $fwrite(32'h80000002,"\n"); // @[LoopBlock.scala 955:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [4:0]  io_InLiveIn_0_bits_taskID,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [4:0]  io_InLiveIn_2_bits_taskID,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [4:0]  io_InLiveIn_3_bits_taskID,
  input  [31:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [4:0]  io_InLiveIn_4_bits_taskID,
  input  [31:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input  [31:0] io_InLiveIn_5_bits_data,
  output        io_InLiveIn_6_ready,
  input         io_InLiveIn_6_valid,
  input  [4:0]  io_InLiveIn_6_bits_taskID,
  input  [31:0] io_InLiveIn_6_bits_data,
  output        io_InLiveIn_7_ready,
  input         io_InLiveIn_7_valid,
  input  [31:0] io_InLiveIn_7_bits_data,
  output        io_InLiveIn_8_ready,
  input         io_InLiveIn_8_valid,
  input  [4:0]  io_InLiveIn_8_bits_taskID,
  input  [31:0] io_InLiveIn_8_bits_data,
  output        io_InLiveIn_9_ready,
  input         io_InLiveIn_9_valid,
  input  [31:0] io_InLiveIn_9_bits_data,
  output        io_InLiveIn_10_ready,
  input         io_InLiveIn_10_valid,
  input  [31:0] io_InLiveIn_10_bits_data,
  output        io_InLiveIn_11_ready,
  input         io_InLiveIn_11_valid,
  input  [4:0]  io_InLiveIn_11_bits_taskID,
  input  [31:0] io_InLiveIn_11_bits_data,
  output        io_InLiveIn_12_ready,
  input         io_InLiveIn_12_valid,
  input  [31:0] io_InLiveIn_12_bits_data,
  output        io_InLiveIn_13_ready,
  input         io_InLiveIn_13_valid,
  input  [31:0] io_InLiveIn_13_bits_data,
  output        io_InLiveIn_14_ready,
  input         io_InLiveIn_14_valid,
  input  [31:0] io_InLiveIn_14_bits_data,
  input         io_OutLiveIn_field14_0_ready,
  output        io_OutLiveIn_field14_0_valid,
  output [31:0] io_OutLiveIn_field14_0_bits_data,
  input         io_OutLiveIn_field13_0_ready,
  output        io_OutLiveIn_field13_0_valid,
  output [31:0] io_OutLiveIn_field13_0_bits_data,
  input         io_OutLiveIn_field12_0_ready,
  output        io_OutLiveIn_field12_0_valid,
  output [31:0] io_OutLiveIn_field12_0_bits_data,
  input         io_OutLiveIn_field11_0_ready,
  output        io_OutLiveIn_field11_0_valid,
  output [4:0]  io_OutLiveIn_field11_0_bits_taskID,
  output [31:0] io_OutLiveIn_field11_0_bits_data,
  input         io_OutLiveIn_field10_0_ready,
  output        io_OutLiveIn_field10_0_valid,
  output [31:0] io_OutLiveIn_field10_0_bits_data,
  input         io_OutLiveIn_field9_0_ready,
  output        io_OutLiveIn_field9_0_valid,
  output [31:0] io_OutLiveIn_field9_0_bits_data,
  input         io_OutLiveIn_field8_0_ready,
  output        io_OutLiveIn_field8_0_valid,
  output [4:0]  io_OutLiveIn_field8_0_bits_taskID,
  output [31:0] io_OutLiveIn_field8_0_bits_data,
  input         io_OutLiveIn_field7_0_ready,
  output        io_OutLiveIn_field7_0_valid,
  output [31:0] io_OutLiveIn_field7_0_bits_data,
  input         io_OutLiveIn_field6_0_ready,
  output        io_OutLiveIn_field6_0_valid,
  output [4:0]  io_OutLiveIn_field6_0_bits_taskID,
  output [31:0] io_OutLiveIn_field6_0_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output [31:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [4:0]  io_OutLiveIn_field4_0_bits_taskID,
  output [31:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [4:0]  io_OutLiveIn_field3_0_bits_taskID,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [4:0]  io_OutLiveIn_field2_0_bits_taskID,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [4:0]  io_OutLiveIn_field0_0_bits_taskID,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_OutLiveIn_field0_1_ready,
  output        io_OutLiveIn_field0_1_valid,
  output [31:0] io_OutLiveIn_field0_1_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_2;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_3;
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_5;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_6;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_7;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_8;
  reg [4:0] in_live_in_R_0_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [4:0] in_live_in_R_2_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [4:0] in_live_in_R_3_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_15;
  reg [4:0] in_live_in_R_4_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_16;
  reg [31:0] in_live_in_R_4_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_17;
  reg [31:0] in_live_in_R_5_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_18;
  reg [4:0] in_live_in_R_6_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_19;
  reg [31:0] in_live_in_R_6_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_20;
  reg [31:0] in_live_in_R_7_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_21;
  reg [4:0] in_live_in_R_8_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_22;
  reg [31:0] in_live_in_R_8_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_23;
  reg [31:0] in_live_in_R_9_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_24;
  reg [31:0] in_live_in_R_10_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_25;
  reg [4:0] in_live_in_R_11_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_26;
  reg [31:0] in_live_in_R_11_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_27;
  reg [31:0] in_live_in_R_12_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_28;
  reg [31:0] in_live_in_R_13_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_29;
  reg [31:0] in_live_in_R_14_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_30;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_31;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_32;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_33;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_34;
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_35;
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_36;
  reg  in_live_in_valid_R_6; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_37;
  reg  in_live_in_valid_R_7; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_38;
  reg  in_live_in_valid_R_8; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_39;
  reg  in_live_in_valid_R_9; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_40;
  reg  in_live_in_valid_R_10; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_41;
  reg  in_live_in_valid_R_11; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_42;
  reg  in_live_in_valid_R_12; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_43;
  reg  in_live_in_valid_R_13; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_44;
  reg  in_live_in_valid_R_14; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_45;
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_46;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_47;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_48;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_49;
  reg  out_live_in_valid_R_0_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_50;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_51;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_52;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_53;
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_54;
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_55;
  reg  out_live_in_valid_R_6_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_56;
  reg  out_live_in_valid_R_7_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_57;
  reg  out_live_in_valid_R_8_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_58;
  reg  out_live_in_valid_R_9_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_59;
  reg  out_live_in_valid_R_10_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_60;
  reg  out_live_in_valid_R_11_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_61;
  reg  out_live_in_valid_R_12_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_62;
  reg  out_live_in_valid_R_13_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_63;
  reg  out_live_in_valid_R_14_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_64;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_65;
  reg  out_live_in_fire_R_0_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_66;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_67;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_68;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_69;
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_70;
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_71;
  reg  out_live_in_fire_R_6_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_72;
  reg  out_live_in_fire_R_7_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_73;
  reg  out_live_in_fire_R_8_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_74;
  reg  out_live_in_fire_R_9_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_75;
  reg  out_live_in_fire_R_10_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_76;
  reg  out_live_in_fire_R_11_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_77;
  reg  out_live_in_fire_R_12_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_78;
  reg  out_live_in_fire_R_13_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_79;
  reg  out_live_in_fire_R_14_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_80;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_81;
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_82;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_83;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_84;
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_85;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_86;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_87;
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_88;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_89;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_90;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_91;
  wire  _T_27; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_29; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[LoopBlock.scala 603:33]
  wire [4:0] _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_31; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_33; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_35; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_37; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_39; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_41; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[LoopBlock.scala 623:33]
  wire  _T_43; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[LoopBlock.scala 623:33]
  wire  _T_45; // @[Decoupled.scala 40:37]
  wire  _GEN_37; // @[LoopBlock.scala 623:33]
  wire  _T_47; // @[Decoupled.scala 40:37]
  wire  _GEN_41; // @[LoopBlock.scala 623:33]
  wire  _T_49; // @[Decoupled.scala 40:37]
  wire  _GEN_45; // @[LoopBlock.scala 623:33]
  wire  _T_51; // @[Decoupled.scala 40:37]
  wire  _GEN_49; // @[LoopBlock.scala 623:33]
  wire  _T_53; // @[Decoupled.scala 40:37]
  wire  _GEN_53; // @[LoopBlock.scala 623:33]
  wire  _T_55; // @[Decoupled.scala 40:37]
  wire  _GEN_57; // @[LoopBlock.scala 623:33]
  wire  _T_57; // @[Decoupled.scala 40:37]
  wire  _GEN_61; // @[LoopBlock.scala 623:33]
  wire  _T_59; // @[Decoupled.scala 40:37]
  wire  _GEN_65; // @[LoopBlock.scala 623:33]
  wire  _T_61; // @[Decoupled.scala 40:37]
  wire  _GEN_69; // @[LoopBlock.scala 623:33]
  wire  _T_63; // @[Decoupled.scala 40:37]
  wire  _GEN_73; // @[LoopBlock.scala 641:37]
  wire  _T_64; // @[Decoupled.scala 40:37]
  wire  _GEN_74; // @[LoopBlock.scala 704:39]
  wire  _T_65; // @[Decoupled.scala 40:37]
  wire  _GEN_75; // @[LoopBlock.scala 708:38]
  wire  _T_66; // @[Decoupled.scala 40:37]
  wire  _GEN_76; // @[LoopBlock.scala 713:33]
  wire  _GEN_77; // @[LoopBlock.scala 713:33]
  wire  _T_67; // @[Decoupled.scala 40:37]
  wire  _GEN_78; // @[LoopBlock.scala 722:57]
  wire  _GEN_79; // @[LoopBlock.scala 722:57]
  wire  _T_68; // @[Decoupled.scala 40:37]
  wire  _GEN_80; // @[LoopBlock.scala 722:57]
  wire  _GEN_81; // @[LoopBlock.scala 722:57]
  wire  _T_69; // @[Decoupled.scala 40:37]
  wire  _GEN_82; // @[LoopBlock.scala 722:57]
  wire  _GEN_83; // @[LoopBlock.scala 722:57]
  wire  _T_70; // @[Decoupled.scala 40:37]
  wire  _GEN_84; // @[LoopBlock.scala 722:57]
  wire  _GEN_85; // @[LoopBlock.scala 722:57]
  wire  _T_71; // @[Decoupled.scala 40:37]
  wire  _GEN_86; // @[LoopBlock.scala 722:57]
  wire  _GEN_87; // @[LoopBlock.scala 722:57]
  wire  _T_72; // @[Decoupled.scala 40:37]
  wire  _GEN_88; // @[LoopBlock.scala 722:57]
  wire  _GEN_89; // @[LoopBlock.scala 722:57]
  wire  _T_73; // @[Decoupled.scala 40:37]
  wire  _GEN_90; // @[LoopBlock.scala 722:57]
  wire  _GEN_91; // @[LoopBlock.scala 722:57]
  wire  _T_74; // @[Decoupled.scala 40:37]
  wire  _GEN_92; // @[LoopBlock.scala 722:57]
  wire  _GEN_93; // @[LoopBlock.scala 722:57]
  wire  _T_75; // @[Decoupled.scala 40:37]
  wire  _GEN_94; // @[LoopBlock.scala 722:57]
  wire  _GEN_95; // @[LoopBlock.scala 722:57]
  wire  _T_76; // @[Decoupled.scala 40:37]
  wire  _GEN_96; // @[LoopBlock.scala 722:57]
  wire  _GEN_97; // @[LoopBlock.scala 722:57]
  wire  _T_77; // @[Decoupled.scala 40:37]
  wire  _GEN_98; // @[LoopBlock.scala 722:57]
  wire  _GEN_99; // @[LoopBlock.scala 722:57]
  wire  _T_78; // @[Decoupled.scala 40:37]
  wire  _GEN_100; // @[LoopBlock.scala 722:57]
  wire  _GEN_101; // @[LoopBlock.scala 722:57]
  wire  _T_79; // @[Decoupled.scala 40:37]
  wire  _GEN_102; // @[LoopBlock.scala 722:57]
  wire  _GEN_103; // @[LoopBlock.scala 722:57]
  wire  _T_80; // @[Decoupled.scala 40:37]
  wire  _GEN_104; // @[LoopBlock.scala 722:57]
  wire  _GEN_105; // @[LoopBlock.scala 722:57]
  wire  _T_81; // @[Decoupled.scala 40:37]
  wire  _GEN_106; // @[LoopBlock.scala 722:57]
  wire  _GEN_107; // @[LoopBlock.scala 722:57]
  wire  _T_82; // @[Decoupled.scala 40:37]
  wire  _GEN_108; // @[LoopBlock.scala 722:57]
  wire  _GEN_109; // @[LoopBlock.scala 722:57]
  wire  _T_83; // @[Decoupled.scala 40:37]
  wire  _GEN_110; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_92;
  wire  _T_84; // @[Conditional.scala 37:30]
  wire  _T_85; // @[LoopBlock.scala 765:35]
  wire  _T_86; // @[LoopBlock.scala 765:35]
  wire  _T_87; // @[LoopBlock.scala 765:35]
  wire  _T_88; // @[LoopBlock.scala 765:35]
  wire  _T_89; // @[LoopBlock.scala 765:35]
  wire  _T_90; // @[LoopBlock.scala 765:35]
  wire  _T_91; // @[LoopBlock.scala 765:35]
  wire  _T_92; // @[LoopBlock.scala 765:35]
  wire  _T_93; // @[LoopBlock.scala 765:35]
  wire  _T_94; // @[LoopBlock.scala 765:35]
  wire  _T_95; // @[LoopBlock.scala 765:35]
  wire  _T_96; // @[LoopBlock.scala 765:35]
  wire  _T_97; // @[LoopBlock.scala 765:35]
  wire  _T_98; // @[LoopBlock.scala 765:35]
  wire  _T_99; // @[LoopBlock.scala 869:28]
  wire  _GEN_112; // @[LoopBlock.scala 870:26]
  wire  _GEN_113; // @[LoopBlock.scala 870:26]
  wire  _GEN_114; // @[LoopBlock.scala 870:26]
  wire  _GEN_115; // @[LoopBlock.scala 870:26]
  wire  _GEN_116; // @[LoopBlock.scala 870:26]
  wire  _GEN_117; // @[LoopBlock.scala 870:26]
  wire  _GEN_118; // @[LoopBlock.scala 870:26]
  wire  _GEN_119; // @[LoopBlock.scala 870:26]
  wire  _GEN_120; // @[LoopBlock.scala 870:26]
  wire  _GEN_121; // @[LoopBlock.scala 870:26]
  wire  _GEN_122; // @[LoopBlock.scala 870:26]
  wire  _GEN_123; // @[LoopBlock.scala 870:26]
  wire  _GEN_124; // @[LoopBlock.scala 870:26]
  wire  _GEN_125; // @[LoopBlock.scala 870:26]
  wire  _GEN_126; // @[LoopBlock.scala 870:26]
  wire  _GEN_127; // @[LoopBlock.scala 870:26]
  wire  _GEN_128; // @[LoopBlock.scala 870:26]
  wire  _GEN_129; // @[LoopBlock.scala 870:26]
  wire  _GEN_131; // @[LoopBlock.scala 870:26]
  wire  _GEN_134; // @[LoopBlock.scala 870:26]
  wire  _GEN_136; // @[LoopBlock.scala 870:26]
  wire  _T_103; // @[Conditional.scala 37:30]
  wire  _T_104; // @[LoopBlock.scala 898:30]
  wire  _T_106; // @[LoopBlock.scala 825:65]
  wire  _T_107; // @[LoopBlock.scala 828:26]
  wire  _T_108; // @[LoopBlock.scala 828:26]
  wire  _T_109; // @[LoopBlock.scala 828:26]
  wire  _T_110; // @[LoopBlock.scala 828:26]
  wire  _T_111; // @[LoopBlock.scala 828:26]
  wire  _T_112; // @[LoopBlock.scala 828:26]
  wire  _T_113; // @[LoopBlock.scala 828:26]
  wire  _T_114; // @[LoopBlock.scala 828:26]
  wire  _T_115; // @[LoopBlock.scala 828:26]
  wire  _T_116; // @[LoopBlock.scala 828:26]
  wire  _T_117; // @[LoopBlock.scala 828:26]
  wire  _T_118; // @[LoopBlock.scala 828:26]
  wire  _T_119; // @[LoopBlock.scala 828:26]
  wire  _T_120; // @[LoopBlock.scala 828:26]
  wire  _T_121; // @[LoopBlock.scala 899:29]
  wire  _T_128; // @[LoopBlock.scala 932:19]
  wire  _T_129; // @[LoopBlock.scala 932:19]
  wire  _GEN_166; // @[LoopBlock.scala 936:64]
  wire  _GEN_169; // @[LoopBlock.scala 936:64]
  wire  _GEN_171; // @[LoopBlock.scala 936:64]
  wire  _GEN_176; // @[LoopBlock.scala 903:56]
  wire  _GEN_177; // @[LoopBlock.scala 903:56]
  wire  _GEN_179; // @[LoopBlock.scala 903:56]
  wire  _GEN_197; // @[LoopBlock.scala 903:56]
  wire  _GEN_198; // @[LoopBlock.scala 903:56]
  wire  _GEN_199; // @[LoopBlock.scala 903:56]
  wire  _GEN_200; // @[LoopBlock.scala 903:56]
  wire  _GEN_201; // @[LoopBlock.scala 903:56]
  wire  _GEN_202; // @[LoopBlock.scala 903:56]
  wire  _GEN_203; // @[LoopBlock.scala 903:56]
  wire  _GEN_204; // @[LoopBlock.scala 903:56]
  wire  _GEN_205; // @[LoopBlock.scala 903:56]
  wire  _GEN_206; // @[LoopBlock.scala 903:56]
  wire  _GEN_207; // @[LoopBlock.scala 903:56]
  wire  _GEN_208; // @[LoopBlock.scala 903:56]
  wire  _GEN_209; // @[LoopBlock.scala 903:56]
  wire  _GEN_210; // @[LoopBlock.scala 903:56]
  wire  _GEN_211; // @[LoopBlock.scala 903:56]
  wire  _GEN_212; // @[LoopBlock.scala 903:56]
  wire  _GEN_213; // @[LoopBlock.scala 903:56]
  wire  _T_137; // @[Conditional.scala 37:30]
  wire  _GEN_646; // @[LoopBlock.scala 932:19]
  wire  _GEN_647; // @[LoopBlock.scala 932:19]
  wire  _GEN_648; // @[LoopBlock.scala 932:19]
  wire  _GEN_649; // @[LoopBlock.scala 932:19]
  wire  _GEN_653; // @[LoopBlock.scala 950:19]
  wire  _GEN_654; // @[LoopBlock.scala 950:19]
  wire  _GEN_655; // @[LoopBlock.scala 950:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_27 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_27 | enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_29 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_29 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_29 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_29 | loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_31 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_31 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_31 | loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_33 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_33 | in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_35 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_35 | in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_37 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_37 | in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_39 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_39 | in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_41 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_41 | in_live_in_valid_R_4; // @[LoopBlock.scala 623:33]
  assign _T_43 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_43 | in_live_in_valid_R_5; // @[LoopBlock.scala 623:33]
  assign _T_45 = io_InLiveIn_6_ready & io_InLiveIn_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_37 = _T_45 | in_live_in_valid_R_6; // @[LoopBlock.scala 623:33]
  assign _T_47 = io_InLiveIn_7_ready & io_InLiveIn_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_41 = _T_47 | in_live_in_valid_R_7; // @[LoopBlock.scala 623:33]
  assign _T_49 = io_InLiveIn_8_ready & io_InLiveIn_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_45 = _T_49 | in_live_in_valid_R_8; // @[LoopBlock.scala 623:33]
  assign _T_51 = io_InLiveIn_9_ready & io_InLiveIn_9_valid; // @[Decoupled.scala 40:37]
  assign _GEN_49 = _T_51 | in_live_in_valid_R_9; // @[LoopBlock.scala 623:33]
  assign _T_53 = io_InLiveIn_10_ready & io_InLiveIn_10_valid; // @[Decoupled.scala 40:37]
  assign _GEN_53 = _T_53 | in_live_in_valid_R_10; // @[LoopBlock.scala 623:33]
  assign _T_55 = io_InLiveIn_11_ready & io_InLiveIn_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_57 = _T_55 | in_live_in_valid_R_11; // @[LoopBlock.scala 623:33]
  assign _T_57 = io_InLiveIn_12_ready & io_InLiveIn_12_valid; // @[Decoupled.scala 40:37]
  assign _GEN_61 = _T_57 | in_live_in_valid_R_12; // @[LoopBlock.scala 623:33]
  assign _T_59 = io_InLiveIn_13_ready & io_InLiveIn_13_valid; // @[Decoupled.scala 40:37]
  assign _GEN_65 = _T_59 | in_live_in_valid_R_13; // @[LoopBlock.scala 623:33]
  assign _T_61 = io_InLiveIn_14_ready & io_InLiveIn_14_valid; // @[Decoupled.scala 40:37]
  assign _GEN_69 = _T_61 | in_live_in_valid_R_14; // @[LoopBlock.scala 623:33]
  assign _T_63 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_73 = _T_63 | in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_64 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  assign _GEN_74 = _T_64 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_65 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  assign _GEN_75 = _T_65 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_66 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_76 = _T_66 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_77 = _T_66 | loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_67 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_78 = _T_67 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_79 = _T_67 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_68 = io_OutLiveIn_field0_1_ready & io_OutLiveIn_field0_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_80 = _T_68 ? 1'h0 : out_live_in_valid_R_0_1; // @[LoopBlock.scala 722:57]
  assign _GEN_81 = _T_68 | out_live_in_fire_R_0_1; // @[LoopBlock.scala 722:57]
  assign _T_69 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_82 = _T_69 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_83 = _T_69 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_70 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_84 = _T_70 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_85 = _T_70 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_71 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_86 = _T_71 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_87 = _T_71 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_72 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_88 = _T_72 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 722:57]
  assign _GEN_89 = _T_72 | out_live_in_fire_R_4_0; // @[LoopBlock.scala 722:57]
  assign _T_73 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_90 = _T_73 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 722:57]
  assign _GEN_91 = _T_73 | out_live_in_fire_R_5_0; // @[LoopBlock.scala 722:57]
  assign _T_74 = io_OutLiveIn_field6_0_ready & io_OutLiveIn_field6_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_92 = _T_74 ? 1'h0 : out_live_in_valid_R_6_0; // @[LoopBlock.scala 722:57]
  assign _GEN_93 = _T_74 | out_live_in_fire_R_6_0; // @[LoopBlock.scala 722:57]
  assign _T_75 = io_OutLiveIn_field7_0_ready & io_OutLiveIn_field7_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_94 = _T_75 ? 1'h0 : out_live_in_valid_R_7_0; // @[LoopBlock.scala 722:57]
  assign _GEN_95 = _T_75 | out_live_in_fire_R_7_0; // @[LoopBlock.scala 722:57]
  assign _T_76 = io_OutLiveIn_field8_0_ready & io_OutLiveIn_field8_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_96 = _T_76 ? 1'h0 : out_live_in_valid_R_8_0; // @[LoopBlock.scala 722:57]
  assign _GEN_97 = _T_76 | out_live_in_fire_R_8_0; // @[LoopBlock.scala 722:57]
  assign _T_77 = io_OutLiveIn_field9_0_ready & io_OutLiveIn_field9_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_98 = _T_77 ? 1'h0 : out_live_in_valid_R_9_0; // @[LoopBlock.scala 722:57]
  assign _GEN_99 = _T_77 | out_live_in_fire_R_9_0; // @[LoopBlock.scala 722:57]
  assign _T_78 = io_OutLiveIn_field10_0_ready & io_OutLiveIn_field10_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_100 = _T_78 ? 1'h0 : out_live_in_valid_R_10_0; // @[LoopBlock.scala 722:57]
  assign _GEN_101 = _T_78 | out_live_in_fire_R_10_0; // @[LoopBlock.scala 722:57]
  assign _T_79 = io_OutLiveIn_field11_0_ready & io_OutLiveIn_field11_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_102 = _T_79 ? 1'h0 : out_live_in_valid_R_11_0; // @[LoopBlock.scala 722:57]
  assign _GEN_103 = _T_79 | out_live_in_fire_R_11_0; // @[LoopBlock.scala 722:57]
  assign _T_80 = io_OutLiveIn_field12_0_ready & io_OutLiveIn_field12_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_104 = _T_80 ? 1'h0 : out_live_in_valid_R_12_0; // @[LoopBlock.scala 722:57]
  assign _GEN_105 = _T_80 | out_live_in_fire_R_12_0; // @[LoopBlock.scala 722:57]
  assign _T_81 = io_OutLiveIn_field13_0_ready & io_OutLiveIn_field13_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_106 = _T_81 ? 1'h0 : out_live_in_valid_R_13_0; // @[LoopBlock.scala 722:57]
  assign _GEN_107 = _T_81 | out_live_in_fire_R_13_0; // @[LoopBlock.scala 722:57]
  assign _T_82 = io_OutLiveIn_field14_0_ready & io_OutLiveIn_field14_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_108 = _T_82 ? 1'h0 : out_live_in_valid_R_14_0; // @[LoopBlock.scala 722:57]
  assign _GEN_109 = _T_82 | out_live_in_fire_R_14_0; // @[LoopBlock.scala 722:57]
  assign _T_83 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_110 = _T_83 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_84 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_85 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_86 = _T_85 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_87 = _T_86 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_88 = _T_87 & in_live_in_valid_R_4; // @[LoopBlock.scala 765:35]
  assign _T_89 = _T_88 & in_live_in_valid_R_5; // @[LoopBlock.scala 765:35]
  assign _T_90 = _T_89 & in_live_in_valid_R_6; // @[LoopBlock.scala 765:35]
  assign _T_91 = _T_90 & in_live_in_valid_R_7; // @[LoopBlock.scala 765:35]
  assign _T_92 = _T_91 & in_live_in_valid_R_8; // @[LoopBlock.scala 765:35]
  assign _T_93 = _T_92 & in_live_in_valid_R_9; // @[LoopBlock.scala 765:35]
  assign _T_94 = _T_93 & in_live_in_valid_R_10; // @[LoopBlock.scala 765:35]
  assign _T_95 = _T_94 & in_live_in_valid_R_11; // @[LoopBlock.scala 765:35]
  assign _T_96 = _T_95 & in_live_in_valid_R_12; // @[LoopBlock.scala 765:35]
  assign _T_97 = _T_96 & in_live_in_valid_R_13; // @[LoopBlock.scala 765:35]
  assign _T_98 = _T_97 & in_live_in_valid_R_14; // @[LoopBlock.scala 765:35]
  assign _T_99 = _T_98 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_112 = enable_R_control | _GEN_78; // @[LoopBlock.scala 870:26]
  assign _GEN_113 = enable_R_control | _GEN_80; // @[LoopBlock.scala 870:26]
  assign _GEN_114 = enable_R_control | _GEN_82; // @[LoopBlock.scala 870:26]
  assign _GEN_115 = enable_R_control | _GEN_84; // @[LoopBlock.scala 870:26]
  assign _GEN_116 = enable_R_control | _GEN_86; // @[LoopBlock.scala 870:26]
  assign _GEN_117 = enable_R_control | _GEN_88; // @[LoopBlock.scala 870:26]
  assign _GEN_118 = enable_R_control | _GEN_90; // @[LoopBlock.scala 870:26]
  assign _GEN_119 = enable_R_control | _GEN_92; // @[LoopBlock.scala 870:26]
  assign _GEN_120 = enable_R_control | _GEN_94; // @[LoopBlock.scala 870:26]
  assign _GEN_121 = enable_R_control | _GEN_96; // @[LoopBlock.scala 870:26]
  assign _GEN_122 = enable_R_control | _GEN_98; // @[LoopBlock.scala 870:26]
  assign _GEN_123 = enable_R_control | _GEN_100; // @[LoopBlock.scala 870:26]
  assign _GEN_124 = enable_R_control | _GEN_102; // @[LoopBlock.scala 870:26]
  assign _GEN_125 = enable_R_control | _GEN_104; // @[LoopBlock.scala 870:26]
  assign _GEN_126 = enable_R_control | _GEN_106; // @[LoopBlock.scala 870:26]
  assign _GEN_127 = enable_R_control | _GEN_108; // @[LoopBlock.scala 870:26]
  assign _GEN_128 = enable_R_control | _GEN_110; // @[LoopBlock.scala 870:26]
  assign _GEN_129 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_131 = enable_R_control | _GEN_74; // @[LoopBlock.scala 870:26]
  assign _GEN_134 = enable_R_control | _GEN_75; // @[LoopBlock.scala 870:26]
  assign _GEN_136 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 870:26]
  assign _T_103 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_104 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_106 = out_live_in_fire_R_0_0 & out_live_in_fire_R_0_1; // @[LoopBlock.scala 825:65]
  assign _T_107 = _T_106 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_108 = _T_107 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_109 = _T_108 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_110 = _T_109 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 828:26]
  assign _T_111 = _T_110 & out_live_in_fire_R_5_0; // @[LoopBlock.scala 828:26]
  assign _T_112 = _T_111 & out_live_in_fire_R_6_0; // @[LoopBlock.scala 828:26]
  assign _T_113 = _T_112 & out_live_in_fire_R_7_0; // @[LoopBlock.scala 828:26]
  assign _T_114 = _T_113 & out_live_in_fire_R_8_0; // @[LoopBlock.scala 828:26]
  assign _T_115 = _T_114 & out_live_in_fire_R_9_0; // @[LoopBlock.scala 828:26]
  assign _T_116 = _T_115 & out_live_in_fire_R_10_0; // @[LoopBlock.scala 828:26]
  assign _T_117 = _T_116 & out_live_in_fire_R_11_0; // @[LoopBlock.scala 828:26]
  assign _T_118 = _T_117 & out_live_in_fire_R_12_0; // @[LoopBlock.scala 828:26]
  assign _T_119 = _T_118 & out_live_in_fire_R_13_0; // @[LoopBlock.scala 828:26]
  assign _T_120 = _T_119 & out_live_in_fire_R_14_0; // @[LoopBlock.scala 828:26]
  assign _T_121 = _T_104 & _T_120; // @[LoopBlock.scala 899:29]
  assign _T_128 = $unsigned(reset); // @[LoopBlock.scala 932:19]
  assign _T_129 = _T_128 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_166 = loop_finish_R_0_control | _GEN_76; // @[LoopBlock.scala 936:64]
  assign _GEN_169 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_171 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_176 = loop_back_R_0_control | _GEN_74; // @[LoopBlock.scala 903:56]
  assign _GEN_177 = loop_back_R_0_control | _GEN_169; // @[LoopBlock.scala 903:56]
  assign _GEN_179 = loop_back_R_0_control | _GEN_75; // @[LoopBlock.scala 903:56]
  assign _GEN_197 = loop_back_R_0_control | _GEN_78; // @[LoopBlock.scala 903:56]
  assign _GEN_198 = loop_back_R_0_control | _GEN_80; // @[LoopBlock.scala 903:56]
  assign _GEN_199 = loop_back_R_0_control | _GEN_82; // @[LoopBlock.scala 903:56]
  assign _GEN_200 = loop_back_R_0_control | _GEN_84; // @[LoopBlock.scala 903:56]
  assign _GEN_201 = loop_back_R_0_control | _GEN_86; // @[LoopBlock.scala 903:56]
  assign _GEN_202 = loop_back_R_0_control | _GEN_88; // @[LoopBlock.scala 903:56]
  assign _GEN_203 = loop_back_R_0_control | _GEN_90; // @[LoopBlock.scala 903:56]
  assign _GEN_204 = loop_back_R_0_control | _GEN_92; // @[LoopBlock.scala 903:56]
  assign _GEN_205 = loop_back_R_0_control | _GEN_94; // @[LoopBlock.scala 903:56]
  assign _GEN_206 = loop_back_R_0_control | _GEN_96; // @[LoopBlock.scala 903:56]
  assign _GEN_207 = loop_back_R_0_control | _GEN_98; // @[LoopBlock.scala 903:56]
  assign _GEN_208 = loop_back_R_0_control | _GEN_100; // @[LoopBlock.scala 903:56]
  assign _GEN_209 = loop_back_R_0_control | _GEN_102; // @[LoopBlock.scala 903:56]
  assign _GEN_210 = loop_back_R_0_control | _GEN_104; // @[LoopBlock.scala 903:56]
  assign _GEN_211 = loop_back_R_0_control | _GEN_106; // @[LoopBlock.scala 903:56]
  assign _GEN_212 = loop_back_R_0_control | _GEN_108; // @[LoopBlock.scala 903:56]
  assign _GEN_213 = loop_back_R_0_control | _GEN_110; // @[LoopBlock.scala 903:56]
  assign _T_137 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_4_ready = ~ in_live_in_valid_R_4; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_5_ready = ~ in_live_in_valid_R_5; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_6_ready = ~ in_live_in_valid_R_6; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_7_ready = ~ in_live_in_valid_R_7; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_8_ready = ~ in_live_in_valid_R_8; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_9_ready = ~ in_live_in_valid_R_9; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_10_ready = ~ in_live_in_valid_R_10; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_11_ready = ~ in_live_in_valid_R_11; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_12_ready = ~ in_live_in_valid_R_12; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_13_ready = ~ in_live_in_valid_R_13; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_14_ready = ~ in_live_in_valid_R_14; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field14_0_valid = out_live_in_valid_R_14_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field14_0_bits_data = in_live_in_R_14_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field13_0_valid = out_live_in_valid_R_13_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field13_0_bits_data = in_live_in_R_13_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field12_0_valid = out_live_in_valid_R_12_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field12_0_bits_data = in_live_in_R_12_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field11_0_valid = out_live_in_valid_R_11_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field11_0_bits_taskID = in_live_in_R_11_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field11_0_bits_data = in_live_in_R_11_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_0_valid = out_live_in_valid_R_10_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_0_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field9_0_valid = out_live_in_valid_R_9_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field9_0_bits_data = in_live_in_R_9_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_valid = out_live_in_valid_R_8_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field8_0_bits_taskID = in_live_in_R_8_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_bits_data = in_live_in_R_8_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_valid = out_live_in_valid_R_7_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field7_0_bits_data = in_live_in_R_7_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_valid = out_live_in_valid_R_6_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field6_0_bits_taskID = in_live_in_R_6_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_bits_data = in_live_in_R_6_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_0_bits_taskID = in_live_in_R_4_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_taskID = in_live_in_R_3_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_taskID = in_live_in_R_2_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_taskID = in_live_in_R_0_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_1_valid = out_live_in_valid_R_0_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_1_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
  assign _GEN_646 = _T_84 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_647 = _GEN_646 & _T_103; // @[LoopBlock.scala 932:19]
  assign _GEN_648 = _GEN_647 & _T_121; // @[LoopBlock.scala 932:19]
  assign _GEN_649 = _GEN_648 & loop_back_R_0_control; // @[LoopBlock.scala 932:19]
  assign _GEN_653 = loop_back_R_0_control == 1'h0; // @[LoopBlock.scala 950:19]
  assign _GEN_654 = _GEN_648 & _GEN_653; // @[LoopBlock.scala 950:19]
  assign _GEN_655 = _GEN_654 & loop_finish_R_0_control; // @[LoopBlock.scala 950:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_0_taskID = _RAND_9[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_2_taskID = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_3_taskID = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_R_4_taskID = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_R_4_data = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_R_5_data = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_live_in_R_6_taskID = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_live_in_R_6_data = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_live_in_R_7_data = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_live_in_R_8_taskID = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_live_in_R_8_data = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_live_in_R_9_data = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_live_in_R_10_data = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  in_live_in_R_11_taskID = _RAND_26[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  in_live_in_R_11_data = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  in_live_in_R_12_data = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  in_live_in_R_13_data = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  in_live_in_R_14_data = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  in_live_in_valid_R_6 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  in_live_in_valid_R_7 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  in_live_in_valid_R_8 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  in_live_in_valid_R_9 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  in_live_in_valid_R_10 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  in_live_in_valid_R_11 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  in_live_in_valid_R_12 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  in_live_in_valid_R_13 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  in_live_in_valid_R_14 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_46[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  out_live_in_valid_R_0_1 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  out_live_in_valid_R_6_0 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  out_live_in_valid_R_7_0 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  out_live_in_valid_R_8_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  out_live_in_valid_R_9_0 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  out_live_in_valid_R_10_0 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  out_live_in_valid_R_11_0 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  out_live_in_valid_R_12_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  out_live_in_valid_R_13_0 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  out_live_in_valid_R_14_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  out_live_in_fire_R_0_1 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  out_live_in_fire_R_6_0 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  out_live_in_fire_R_7_0 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  out_live_in_fire_R_8_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  out_live_in_fire_R_9_0 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  out_live_in_fire_R_10_0 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  out_live_in_fire_R_11_0 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  out_live_in_fire_R_12_0 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  out_live_in_fire_R_13_0 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  out_live_in_fire_R_14_0 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_82[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_85[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_88[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  state = _RAND_92[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_27) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_103) begin
          if (_T_27) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_27) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_27) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_27) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_103) begin
          if (_T_27) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_27) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_27) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_84) begin
        enable_valid_R <= _GEN_3;
      end else begin
        if (_T_103) begin
          enable_valid_R <= _GEN_3;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_3;
            end
          end else begin
            enable_valid_R <= _GEN_3;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_29) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_29) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_29) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_29) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_29) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_29) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_29) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_29) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        loop_back_valid_R_0 <= _GEN_6;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_31) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_31) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_31) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_31) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_7;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        loop_finish_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_33) begin
          in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
        end
      end else begin
        if (_T_103) begin
          if (_T_33) begin
            in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_taskID <= 5'h0;
            end else begin
              if (_T_33) begin
                in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
              end
            end
          end else begin
            if (_T_33) begin
              in_live_in_R_0_taskID <= io_InLiveIn_0_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_33) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_33) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_33) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_33) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_35) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_35) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_35) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_35) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_37) begin
          in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
        end
      end else begin
        if (_T_103) begin
          if (_T_37) begin
            in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_taskID <= 5'h0;
            end else begin
              if (_T_37) begin
                in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
              end
            end
          end else begin
            if (_T_37) begin
              in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_37) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_37) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_37) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_37) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_39) begin
          in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
        end
      end else begin
        if (_T_103) begin
          if (_T_39) begin
            in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_taskID <= 5'h0;
            end else begin
              if (_T_39) begin
                in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
              end
            end
          end else begin
            if (_T_39) begin
              in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_39) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_39) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_39) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_39) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_41) begin
          in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
        end
      end else begin
        if (_T_103) begin
          if (_T_41) begin
            in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_taskID <= 5'h0;
            end else begin
              if (_T_41) begin
                in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
              end
            end
          end else begin
            if (_T_41) begin
              in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_41) begin
          in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_41) begin
            in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_data <= 32'h0;
            end else begin
              if (_T_41) begin
                in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
              end
            end
          end else begin
            if (_T_41) begin
              in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_43) begin
          in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_43) begin
            in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_data <= 32'h0;
            end else begin
              if (_T_43) begin
                in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
              end
            end
          end else begin
            if (_T_43) begin
              in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_45) begin
          in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
        end
      end else begin
        if (_T_103) begin
          if (_T_45) begin
            in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_taskID <= 5'h0;
            end else begin
              if (_T_45) begin
                in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
              end
            end
          end else begin
            if (_T_45) begin
              in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_45) begin
          in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_45) begin
            in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_data <= 32'h0;
            end else begin
              if (_T_45) begin
                in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
              end
            end
          end else begin
            if (_T_45) begin
              in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_47) begin
          in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_47) begin
            in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_data <= 32'h0;
            end else begin
              if (_T_47) begin
                in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
              end
            end
          end else begin
            if (_T_47) begin
              in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_49) begin
          in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
        end
      end else begin
        if (_T_103) begin
          if (_T_49) begin
            in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_taskID <= 5'h0;
            end else begin
              if (_T_49) begin
                in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
              end
            end
          end else begin
            if (_T_49) begin
              in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_49) begin
          in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_49) begin
            in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_data <= 32'h0;
            end else begin
              if (_T_49) begin
                in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
              end
            end
          end else begin
            if (_T_49) begin
              in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_9_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_51) begin
          in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_51) begin
            in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_9_data <= 32'h0;
            end else begin
              if (_T_51) begin
                in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
              end
            end
          end else begin
            if (_T_51) begin
              in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_10_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_53) begin
          in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_53) begin
            in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_10_data <= 32'h0;
            end else begin
              if (_T_53) begin
                in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
              end
            end
          end else begin
            if (_T_53) begin
              in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_11_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_55) begin
          in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
        end
      end else begin
        if (_T_103) begin
          if (_T_55) begin
            in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_11_taskID <= 5'h0;
            end else begin
              if (_T_55) begin
                in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
              end
            end
          end else begin
            if (_T_55) begin
              in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_11_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_55) begin
          in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_55) begin
            in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_11_data <= 32'h0;
            end else begin
              if (_T_55) begin
                in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
              end
            end
          end else begin
            if (_T_55) begin
              in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_12_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_57) begin
          in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_57) begin
            in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_12_data <= 32'h0;
            end else begin
              if (_T_57) begin
                in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
              end
            end
          end else begin
            if (_T_57) begin
              in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_13_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_59) begin
          in_live_in_R_13_data <= io_InLiveIn_13_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_59) begin
            in_live_in_R_13_data <= io_InLiveIn_13_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_13_data <= 32'h0;
            end else begin
              if (_T_59) begin
                in_live_in_R_13_data <= io_InLiveIn_13_bits_data;
              end
            end
          end else begin
            if (_T_59) begin
              in_live_in_R_13_data <= io_InLiveIn_13_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_14_data <= 32'h0;
    end else begin
      if (_T_84) begin
        if (_T_61) begin
          in_live_in_R_14_data <= io_InLiveIn_14_bits_data;
        end
      end else begin
        if (_T_103) begin
          if (_T_61) begin
            in_live_in_R_14_data <= io_InLiveIn_14_bits_data;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_14_data <= 32'h0;
            end else begin
              if (_T_61) begin
                in_live_in_R_14_data <= io_InLiveIn_14_bits_data;
              end
            end
          end else begin
            if (_T_61) begin
              in_live_in_R_14_data <= io_InLiveIn_14_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_0 <= _GEN_13;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_0 <= _GEN_13;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              in_live_in_valid_R_0 <= _GEN_13;
            end
          end else begin
            in_live_in_valid_R_0 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_1 <= _GEN_17;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_1 <= _GEN_17;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              in_live_in_valid_R_1 <= _GEN_17;
            end
          end else begin
            in_live_in_valid_R_1 <= _GEN_17;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_2 <= _GEN_21;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              in_live_in_valid_R_2 <= _GEN_21;
            end
          end else begin
            in_live_in_valid_R_2 <= _GEN_21;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_3 <= _GEN_25;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_3 <= _GEN_25;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              in_live_in_valid_R_3 <= _GEN_25;
            end
          end else begin
            in_live_in_valid_R_3 <= _GEN_25;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_4 <= _GEN_29;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_4 <= _GEN_29;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_4 <= 1'h0;
            end else begin
              in_live_in_valid_R_4 <= _GEN_29;
            end
          end else begin
            in_live_in_valid_R_4 <= _GEN_29;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_5 <= _GEN_33;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_5 <= _GEN_33;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_5 <= 1'h0;
            end else begin
              in_live_in_valid_R_5 <= _GEN_33;
            end
          end else begin
            in_live_in_valid_R_5 <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_6 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_6 <= _GEN_37;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_6 <= _GEN_37;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_6 <= 1'h0;
            end else begin
              in_live_in_valid_R_6 <= _GEN_37;
            end
          end else begin
            in_live_in_valid_R_6 <= _GEN_37;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_7 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_7 <= _GEN_41;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_7 <= _GEN_41;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_7 <= 1'h0;
            end else begin
              in_live_in_valid_R_7 <= _GEN_41;
            end
          end else begin
            in_live_in_valid_R_7 <= _GEN_41;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_8 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_8 <= _GEN_45;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_8 <= _GEN_45;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_8 <= 1'h0;
            end else begin
              in_live_in_valid_R_8 <= _GEN_45;
            end
          end else begin
            in_live_in_valid_R_8 <= _GEN_45;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_9 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_9 <= _GEN_49;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_9 <= _GEN_49;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_9 <= 1'h0;
            end else begin
              in_live_in_valid_R_9 <= _GEN_49;
            end
          end else begin
            in_live_in_valid_R_9 <= _GEN_49;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_10 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_10 <= _GEN_53;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_10 <= _GEN_53;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_10 <= 1'h0;
            end else begin
              in_live_in_valid_R_10 <= _GEN_53;
            end
          end else begin
            in_live_in_valid_R_10 <= _GEN_53;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_11 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_11 <= _GEN_57;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_11 <= _GEN_57;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_11 <= 1'h0;
            end else begin
              in_live_in_valid_R_11 <= _GEN_57;
            end
          end else begin
            in_live_in_valid_R_11 <= _GEN_57;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_12 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_12 <= _GEN_61;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_12 <= _GEN_61;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_12 <= 1'h0;
            end else begin
              in_live_in_valid_R_12 <= _GEN_61;
            end
          end else begin
            in_live_in_valid_R_12 <= _GEN_61;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_13 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_13 <= _GEN_65;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_13 <= _GEN_65;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_13 <= 1'h0;
            end else begin
              in_live_in_valid_R_13 <= _GEN_65;
            end
          end else begin
            in_live_in_valid_R_13 <= _GEN_65;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_14 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_live_in_valid_R_14 <= _GEN_69;
      end else begin
        if (_T_103) begin
          in_live_in_valid_R_14 <= _GEN_69;
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_14 <= 1'h0;
            end else begin
              in_live_in_valid_R_14 <= _GEN_69;
            end
          end else begin
            in_live_in_valid_R_14 <= _GEN_69;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_63) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_63) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        in_carry_in_valid_R_0 <= _GEN_73;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_73;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_73;
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_73;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_73;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_0_0 <= _GEN_112;
        end else begin
          if (_T_67) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_0_0 <= _GEN_197;
          end else begin
            if (_T_67) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_67) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_1 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_0_1 <= _GEN_113;
        end else begin
          if (_T_68) begin
            out_live_in_valid_R_0_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_0_1 <= _GEN_198;
          end else begin
            if (_T_68) begin
              out_live_in_valid_R_0_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_68) begin
            out_live_in_valid_R_0_1 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_1_0 <= _GEN_114;
        end else begin
          if (_T_69) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_1_0 <= _GEN_199;
          end else begin
            if (_T_69) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_69) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_2_0 <= _GEN_115;
        end else begin
          if (_T_70) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_2_0 <= _GEN_200;
          end else begin
            if (_T_70) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_70) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_3_0 <= _GEN_116;
        end else begin
          if (_T_71) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_3_0 <= _GEN_201;
          end else begin
            if (_T_71) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_71) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_4_0 <= _GEN_117;
        end else begin
          if (_T_72) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_4_0 <= _GEN_202;
          end else begin
            if (_T_72) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_72) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_5_0 <= _GEN_118;
        end else begin
          if (_T_73) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_5_0 <= _GEN_203;
          end else begin
            if (_T_73) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_73) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_6_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_6_0 <= _GEN_119;
        end else begin
          if (_T_74) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_6_0 <= _GEN_204;
          end else begin
            if (_T_74) begin
              out_live_in_valid_R_6_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_74) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_7_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_7_0 <= _GEN_120;
        end else begin
          if (_T_75) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_7_0 <= _GEN_205;
          end else begin
            if (_T_75) begin
              out_live_in_valid_R_7_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_75) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_8_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_8_0 <= _GEN_121;
        end else begin
          if (_T_76) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_8_0 <= _GEN_206;
          end else begin
            if (_T_76) begin
              out_live_in_valid_R_8_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_9_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_9_0 <= _GEN_122;
        end else begin
          if (_T_77) begin
            out_live_in_valid_R_9_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_9_0 <= _GEN_207;
          end else begin
            if (_T_77) begin
              out_live_in_valid_R_9_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_77) begin
            out_live_in_valid_R_9_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_10_0 <= _GEN_123;
        end else begin
          if (_T_78) begin
            out_live_in_valid_R_10_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_10_0 <= _GEN_208;
          end else begin
            if (_T_78) begin
              out_live_in_valid_R_10_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_78) begin
            out_live_in_valid_R_10_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_11_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_11_0 <= _GEN_124;
        end else begin
          if (_T_79) begin
            out_live_in_valid_R_11_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_11_0 <= _GEN_209;
          end else begin
            if (_T_79) begin
              out_live_in_valid_R_11_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_79) begin
            out_live_in_valid_R_11_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_12_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_12_0 <= _GEN_125;
        end else begin
          if (_T_80) begin
            out_live_in_valid_R_12_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_12_0 <= _GEN_210;
          end else begin
            if (_T_80) begin
              out_live_in_valid_R_12_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_80) begin
            out_live_in_valid_R_12_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_13_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_13_0 <= _GEN_126;
        end else begin
          if (_T_81) begin
            out_live_in_valid_R_13_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_13_0 <= _GEN_211;
          end else begin
            if (_T_81) begin
              out_live_in_valid_R_13_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_81) begin
            out_live_in_valid_R_13_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_14_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_live_in_valid_R_14_0 <= _GEN_127;
        end else begin
          if (_T_82) begin
            out_live_in_valid_R_14_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_live_in_valid_R_14_0 <= _GEN_212;
          end else begin
            if (_T_82) begin
              out_live_in_valid_R_14_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_82) begin
            out_live_in_valid_R_14_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_0_0 <= _GEN_79;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_0 <= _GEN_79;
            end
          end else begin
            out_live_in_fire_R_0_0 <= _GEN_79;
          end
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_79;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_1 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_0_1 <= _GEN_81;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_1 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_1 <= _GEN_81;
            end
          end else begin
            out_live_in_fire_R_0_1 <= _GEN_81;
          end
        end else begin
          out_live_in_fire_R_0_1 <= _GEN_81;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_1_0 <= _GEN_83;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_0 <= _GEN_83;
            end
          end else begin
            out_live_in_fire_R_1_0 <= _GEN_83;
          end
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_83;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_2_0 <= _GEN_85;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_2_0 <= _GEN_85;
            end
          end else begin
            out_live_in_fire_R_2_0 <= _GEN_85;
          end
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_85;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_3_0 <= _GEN_87;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_3_0 <= _GEN_87;
            end
          end else begin
            out_live_in_fire_R_3_0 <= _GEN_87;
          end
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_87;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_4_0 <= _GEN_89;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_4_0 <= _GEN_89;
            end
          end else begin
            out_live_in_fire_R_4_0 <= _GEN_89;
          end
        end else begin
          out_live_in_fire_R_4_0 <= _GEN_89;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_5_0 <= _GEN_91;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_5_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_5_0 <= _GEN_91;
            end
          end else begin
            out_live_in_fire_R_5_0 <= _GEN_91;
          end
        end else begin
          out_live_in_fire_R_5_0 <= _GEN_91;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_6_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_6_0 <= _GEN_93;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_6_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_6_0 <= _GEN_93;
            end
          end else begin
            out_live_in_fire_R_6_0 <= _GEN_93;
          end
        end else begin
          out_live_in_fire_R_6_0 <= _GEN_93;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_7_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_7_0 <= _GEN_95;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_7_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_7_0 <= _GEN_95;
            end
          end else begin
            out_live_in_fire_R_7_0 <= _GEN_95;
          end
        end else begin
          out_live_in_fire_R_7_0 <= _GEN_95;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_8_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_8_0 <= _GEN_97;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_8_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_8_0 <= _GEN_97;
            end
          end else begin
            out_live_in_fire_R_8_0 <= _GEN_97;
          end
        end else begin
          out_live_in_fire_R_8_0 <= _GEN_97;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_9_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_9_0 <= _GEN_99;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_9_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_9_0 <= _GEN_99;
            end
          end else begin
            out_live_in_fire_R_9_0 <= _GEN_99;
          end
        end else begin
          out_live_in_fire_R_9_0 <= _GEN_99;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_10_0 <= _GEN_101;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_0 <= _GEN_101;
            end
          end else begin
            out_live_in_fire_R_10_0 <= _GEN_101;
          end
        end else begin
          out_live_in_fire_R_10_0 <= _GEN_101;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_11_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_11_0 <= _GEN_103;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_11_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_11_0 <= _GEN_103;
            end
          end else begin
            out_live_in_fire_R_11_0 <= _GEN_103;
          end
        end else begin
          out_live_in_fire_R_11_0 <= _GEN_103;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_12_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_12_0 <= _GEN_105;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_12_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_12_0 <= _GEN_105;
            end
          end else begin
            out_live_in_fire_R_12_0 <= _GEN_105;
          end
        end else begin
          out_live_in_fire_R_12_0 <= _GEN_105;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_13_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_13_0 <= _GEN_107;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_13_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_13_0 <= _GEN_107;
            end
          end else begin
            out_live_in_fire_R_13_0 <= _GEN_107;
          end
        end else begin
          out_live_in_fire_R_13_0 <= _GEN_107;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_14_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        out_live_in_fire_R_14_0 <= _GEN_109;
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_14_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_14_0 <= _GEN_109;
            end
          end else begin
            out_live_in_fire_R_14_0 <= _GEN_109;
          end
        end else begin
          out_live_in_fire_R_14_0 <= _GEN_109;
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          out_carry_out_valid_R_0_0 <= _GEN_128;
        end else begin
          if (_T_83) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            out_carry_out_valid_R_0_0 <= _GEN_213;
          end else begin
            if (_T_83) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_83) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          active_loop_start_R_control <= _GEN_129;
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          active_loop_start_valid_R <= _GEN_131;
        end else begin
          if (_T_64) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            active_loop_start_valid_R <= _GEN_176;
          end else begin
            if (_T_64) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_64) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            active_loop_back_R_control <= _GEN_177;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          active_loop_back_valid_R <= _GEN_134;
        end else begin
          if (_T_65) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            active_loop_back_valid_R <= _GEN_179;
          end else begin
            if (_T_65) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_65) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 5'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          loop_exit_R_0_control <= _GEN_136;
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (!(loop_back_R_0_control)) begin
              loop_exit_R_0_control <= _GEN_171;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          if (enable_R_control) begin
            if (_T_66) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_66) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              if (_T_66) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              loop_exit_valid_R_0 <= _GEN_166;
            end
          end else begin
            if (_T_66) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_76;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_77;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_84) begin
        if (_T_99) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_103) begin
          if (_T_121) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_137) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_649 & _T_129) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_5: Restarted fired @ %d\n",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 932:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_655 & _T_129) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOOP]   Loop_5: Output fired @ %d ",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 950:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_655 & _T_129) begin
          $fwrite(32'h80000002,"\n"); // @[LoopBlock.scala 955:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_valid_R_1; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_6;
  reg  output_valid_R_2; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_7;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_8;
  reg  output_fire_R_1; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_9;
  reg  output_fire_R_2; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_10;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BasicBlock.scala 244:28]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_1; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_2; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_11;
  wire  _T_21; // @[Conditional.scala 37:30]
  wire  _T_25; // @[BasicBlock.scala 309:81]
  wire  _T_26; // @[BasicBlock.scala 309:81]
  wire  _T_27; // @[BasicBlock.scala 309:81]
  wire  _T_28; // @[BasicBlock.scala 315:19]
  wire  _T_29; // @[BasicBlock.scala 315:19]
  wire  _GEN_10; // @[BasicBlock.scala 304:8]
  wire  _GEN_11; // @[BasicBlock.scala 304:8]
  wire  _GEN_12; // @[BasicBlock.scala 304:8]
  wire  _GEN_16; // @[BasicBlock.scala 304:8]
  wire  _T_33; // @[BasicBlock.scala 328:35]
  wire  _T_34; // @[BasicBlock.scala 328:35]
  wire  _GEN_44; // @[BasicBlock.scala 315:19]
  wire  _GEN_45; // @[BasicBlock.scala 315:19]
  wire  _GEN_47; // @[BasicBlock.scala 320:19]
  wire  _GEN_48; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 244:28]
  assign _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 256:85]
  assign _T_21 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_25 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_26 = _T_9 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_27 = _T_10 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_28 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_29 = _T_28 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_10 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_11 = _GEN_3 | output_valid_R_1; // @[BasicBlock.scala 304:8]
  assign _GEN_12 = _GEN_3 | output_valid_R_2; // @[BasicBlock.scala 304:8]
  assign _GEN_16 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign _T_33 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 328:35]
  assign _T_34 = _T_33 & out_fire_mask_2; // @[BasicBlock.scala 328:35]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_21 ? _GEN_10 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_1_valid = _T_21 ? _GEN_11 : output_valid_R_1; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_1_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_2_valid = _T_21 ? _GEN_12 : output_valid_R_2; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_2_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_44 = _T_21 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_45 = _GEN_44 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_47 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_48 = _GEN_44 & _GEN_47; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_21) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_21) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_21) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_34) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_21) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_25;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else begin
      if (_T_21) begin
        if (_GEN_3) begin
          output_valid_R_1 <= _T_26;
        end else begin
          if (_T_9) begin
            output_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_9) begin
          output_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else begin
      if (_T_21) begin
        if (_GEN_3) begin
          output_valid_R_2 <= _T_27;
        end else begin
          if (_T_10) begin
            output_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_10) begin
          output_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_21) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (_T_34) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else begin
      if (_T_21) begin
        output_fire_R_1 <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_34) begin
            output_fire_R_1 <= 1'h0;
          end else begin
            output_fire_R_1 <= _GEN_6;
          end
        end else begin
          output_fire_R_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else begin
      if (_T_21) begin
        output_fire_R_2 <= _GEN_8;
      end else begin
        if (state) begin
          if (_T_34) begin
            output_fire_R_2 <= 1'h0;
          end else begin
            output_fire_R_2 <= _GEN_8;
          end
        end else begin
          output_fire_R_2 <= _GEN_8;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_21) begin
        state <= _GEN_16;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_45 & _T_29) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_entry0: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_48 & _T_29) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_entry0: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_1(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_valid_R_1; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_6;
  reg  output_valid_R_2; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_7;
  reg  output_valid_R_3; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_8;
  reg  output_valid_R_4; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_9;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_10;
  reg  output_fire_R_1; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_11;
  reg  output_fire_R_2; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_12;
  reg  output_fire_R_3; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_13;
  reg  output_fire_R_4; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_14;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BasicBlock.scala 244:28]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[BasicBlock.scala 244:28]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_10; // @[BasicBlock.scala 244:28]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_12; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_1; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_2; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_3; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_4; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_15;
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_33; // @[BasicBlock.scala 309:81]
  wire  _T_34; // @[BasicBlock.scala 309:81]
  wire  _T_35; // @[BasicBlock.scala 309:81]
  wire  _T_36; // @[BasicBlock.scala 309:81]
  wire  _T_37; // @[BasicBlock.scala 309:81]
  wire  _T_38; // @[BasicBlock.scala 315:19]
  wire  _T_39; // @[BasicBlock.scala 315:19]
  wire  _GEN_14; // @[BasicBlock.scala 304:8]
  wire  _GEN_15; // @[BasicBlock.scala 304:8]
  wire  _GEN_16; // @[BasicBlock.scala 304:8]
  wire  _GEN_17; // @[BasicBlock.scala 304:8]
  wire  _GEN_18; // @[BasicBlock.scala 304:8]
  wire  _GEN_24; // @[BasicBlock.scala 304:8]
  wire  _T_43; // @[BasicBlock.scala 328:35]
  wire  _T_44; // @[BasicBlock.scala 328:35]
  wire  _T_45; // @[BasicBlock.scala 328:35]
  wire  _T_46; // @[BasicBlock.scala 328:35]
  wire  _GEN_62; // @[BasicBlock.scala 315:19]
  wire  _GEN_63; // @[BasicBlock.scala 315:19]
  wire  _GEN_65; // @[BasicBlock.scala 320:19]
  wire  _GEN_66; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 244:28]
  assign _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 244:28]
  assign _T_11 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_10 = _T_11 | output_fire_R_3; // @[BasicBlock.scala 244:28]
  assign _T_12 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_12 = _T_12 | output_fire_R_4; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_3 = output_fire_R_3 | _T_11; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_4 = output_fire_R_4 | _T_12; // @[BasicBlock.scala 256:85]
  assign _T_27 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_33 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_34 = _T_9 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_35 = _T_10 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_36 = _T_11 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_37 = _T_12 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_38 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_39 = _T_38 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_14 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_15 = _GEN_3 | output_valid_R_1; // @[BasicBlock.scala 304:8]
  assign _GEN_16 = _GEN_3 | output_valid_R_2; // @[BasicBlock.scala 304:8]
  assign _GEN_17 = _GEN_3 | output_valid_R_3; // @[BasicBlock.scala 304:8]
  assign _GEN_18 = _GEN_3 | output_valid_R_4; // @[BasicBlock.scala 304:8]
  assign _GEN_24 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign _T_43 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 328:35]
  assign _T_44 = _T_43 & out_fire_mask_2; // @[BasicBlock.scala 328:35]
  assign _T_45 = _T_44 & out_fire_mask_3; // @[BasicBlock.scala 328:35]
  assign _T_46 = _T_45 & out_fire_mask_4; // @[BasicBlock.scala 328:35]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_27 ? _GEN_14 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_1_valid = _T_27 ? _GEN_15 : output_valid_R_1; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_1_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_2_valid = _T_27 ? _GEN_16 : output_valid_R_2; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_2_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_3_valid = _T_27 ? _GEN_17 : output_valid_R_3; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_3_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_3_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_4_valid = _T_27 ? _GEN_18 : output_valid_R_4; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_4_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_4_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_62 = _T_27 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_63 = _GEN_62 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_65 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_66 = _GEN_62 & _GEN_65; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_4 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  output_fire_R_4 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_46) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_46) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_27) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_46) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_33;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_1 <= _T_34;
        end else begin
          if (_T_9) begin
            output_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_9) begin
          output_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_2 <= _T_35;
        end else begin
          if (_T_10) begin
            output_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_10) begin
          output_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_3 <= _T_36;
        end else begin
          if (_T_11) begin
            output_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_11) begin
          output_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_4 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_4 <= _T_37;
        end else begin
          if (_T_12) begin
            output_valid_R_4 <= 1'h0;
          end
        end
      end else begin
        if (_T_12) begin
          output_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_1 <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_1 <= 1'h0;
          end else begin
            output_fire_R_1 <= _GEN_6;
          end
        end else begin
          output_fire_R_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_2 <= _GEN_8;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_2 <= 1'h0;
          end else begin
            output_fire_R_2 <= _GEN_8;
          end
        end else begin
          output_fire_R_2 <= _GEN_8;
        end
      end
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_3 <= _GEN_10;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_3 <= 1'h0;
          end else begin
            output_fire_R_3 <= _GEN_10;
          end
        end else begin
          output_fire_R_3 <= _GEN_10;
        end
      end
    end
    if (reset) begin
      output_fire_R_4 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_4 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_4 <= 1'h0;
          end else begin
            output_fire_R_4 <= _GEN_12;
          end
        end else begin
          output_fire_R_4 <= _GEN_12;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_27) begin
        state <= _GEN_24;
      end else begin
        if (state) begin
          if (_T_46) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body_lr_ph1: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body_lr_ph1: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_2(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_6;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_7;
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_17; // @[BasicBlock.scala 309:81]
  wire  _T_18; // @[BasicBlock.scala 315:19]
  wire  _T_19; // @[BasicBlock.scala 315:19]
  wire  _GEN_6; // @[BasicBlock.scala 304:8]
  wire  _GEN_8; // @[BasicBlock.scala 304:8]
  wire  _GEN_26; // @[BasicBlock.scala 315:19]
  wire  _GEN_27; // @[BasicBlock.scala 315:19]
  wire  _GEN_29; // @[BasicBlock.scala 320:19]
  wire  _GEN_30; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_18 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_19 = _T_18 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_6 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_8 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_15 ? _GEN_6 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_26 = _T_15 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_27 = _GEN_26 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_29 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_17;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_8;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup_loopexit2: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup_loopexit2: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_3(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg [4:0] in_data_R_1_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_3;
  reg  in_data_R_1_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_4;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_5;
  reg  in_data_valid_R_1; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_6;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_7;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_8;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_9;
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[BasicBlock.scala 232:36]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 232:36]
  wire  _GEN_6; // @[BasicBlock.scala 232:36]
  wire [4:0] _T_11; // @[BasicBlock.scala 239:34]
  wire [4:0] _T_12; // @[BasicBlock.scala 239:34]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 240:15]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  wire  predicate_val; // @[BasicBlock.scala 264:57]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_10;
  wire  _T_26; // @[Conditional.scala 37:30]
  wire  _T_27; // @[BasicBlock.scala 299:41]
  wire  _T_29; // @[BasicBlock.scala 309:81]
  wire  _T_30; // @[BasicBlock.scala 315:19]
  wire  _T_31; // @[BasicBlock.scala 315:19]
  wire  _GEN_9; // @[BasicBlock.scala 304:8]
  wire  _GEN_11; // @[BasicBlock.scala 304:8]
  wire  _GEN_38; // @[BasicBlock.scala 315:19]
  wire  _GEN_39; // @[BasicBlock.scala 315:19]
  wire  _GEN_41; // @[BasicBlock.scala 320:19]
  wire  _GEN_42; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_8 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_8 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 232:36]
  assign _GEN_3 = _T_8 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign _T_10 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_10 ? io_predicateIn_1_bits_control : in_data_R_1_control; // @[BasicBlock.scala 232:36]
  assign _GEN_6 = _T_10 | in_data_valid_R_1; // @[BasicBlock.scala 232:36]
  assign _T_11 = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_12 = io_predicateIn_1_bits_taskID | in_data_R_1_taskID; // @[BasicBlock.scala 239:34]
  assign in_task_ID = _T_11 | _T_12; // @[BasicBlock.scala 240:15]
  assign _T_13 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_13 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_13; // @[BasicBlock.scala 256:85]
  assign predicate_val = in_data_R_0_control | in_data_R_1_control; // @[BasicBlock.scala 264:57]
  assign _T_26 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_27 = _GEN_3 & _GEN_6; // @[BasicBlock.scala 299:41]
  assign _T_29 = _T_13 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_30 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_31 = _T_30 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_9 = _T_27 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_11 = _T_27 | state; // @[BasicBlock.scala 304:8]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_predicateIn_1_ready = ~ in_data_valid_R_1; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_26 ? _GEN_9 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = _T_11 | _T_12; // @[BasicBlock.scala 282:22]
  assign io_Out_0_bits_control = _GEN_1 | _GEN_4; // @[BasicBlock.scala 282:22]
  assign _GEN_38 = _T_26 & _T_27; // @[BasicBlock.scala 315:19]
  assign _GEN_39 = _GEN_38 & predicate_val; // @[BasicBlock.scala 315:19]
  assign _GEN_41 = predicate_val == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_42 = _GEN_38 & _GEN_41; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_R_1_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_26) begin
        if (_T_8) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_8) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_8) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_26) begin
        if (_T_8) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_8) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_8) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_taskID <= 5'h0;
    end else begin
      if (_T_26) begin
        if (_T_10) begin
          in_data_R_1_taskID <= io_predicateIn_1_bits_taskID;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_1_taskID <= 5'h0;
          end else begin
            if (_T_10) begin
              in_data_R_1_taskID <= io_predicateIn_1_bits_taskID;
            end
          end
        end else begin
          if (_T_10) begin
            in_data_R_1_taskID <= io_predicateIn_1_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_control <= 1'h0;
    end else begin
      if (_T_26) begin
        if (_T_10) begin
          in_data_R_1_control <= io_predicateIn_1_bits_control;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_1_control <= 1'h0;
          end else begin
            if (_T_10) begin
              in_data_R_1_control <= io_predicateIn_1_bits_control;
            end
          end
        end else begin
          if (_T_10) begin
            in_data_R_1_control <= io_predicateIn_1_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_26) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_26) begin
        in_data_valid_R_1 <= _GEN_6;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_6;
          end
        end else begin
          in_data_valid_R_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_26) begin
        if (_T_27) begin
          output_valid_R_0 <= _T_29;
        end else begin
          if (_T_13) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_13) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_26) begin
        output_fire_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_7;
          end
        end else begin
          output_fire_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_26) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_39 & _T_31) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup3: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_31) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup3: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_4;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_5;
  reg  out_valid_R_2; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_6;
  reg  out_valid_R_3; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_7;
  reg  mask_valid_R_0; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_8;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 716:29]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[HandShaking.scala 716:29]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[HandShaking.scala 727:32]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_9;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_10;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_11;
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_12;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_13;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_14;
  reg  predicate_control_R_1; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_15;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_16;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_17;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_18;
  wire  predicate; // @[BasicBlock.scala 75:58]
  wire [4:0] predicate_task; // @[BasicBlock.scala 76:62]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _T_16; // @[BasicBlock.scala 78:91]
  wire  _T_17; // @[BasicBlock.scala 78:91]
  wire  start; // @[BasicBlock.scala 78:107]
  wire [1:0] _T_22; // @[BasicBlock.scala 102:52]
  wire  _T_23; // @[Conditional.scala 37:30]
  wire  _GEN_19; // @[BasicBlock.scala 112:19]
  wire  _GEN_20; // @[BasicBlock.scala 112:19]
  wire  _GEN_21; // @[BasicBlock.scala 112:19]
  wire  _GEN_22; // @[BasicBlock.scala 112:19]
  wire  _GEN_23; // @[BasicBlock.scala 112:19]
  wire  _GEN_24; // @[BasicBlock.scala 112:19]
  wire [3:0] _T_28; // @[HandShaking.scala 741:17]
  wire  _T_29; // @[HandShaking.scala 741:24]
  wire  _T_32; // @[BasicBlock.scala 126:19]
  wire  _T_33; // @[BasicBlock.scala 126:19]
  wire  _GEN_54; // @[BasicBlock.scala 126:19]
  wire  _GEN_55; // @[BasicBlock.scala 126:19]
  wire  _GEN_56; // @[BasicBlock.scala 126:19]
  wire  _GEN_57; // @[BasicBlock.scala 126:19]
  wire  _GEN_61; // @[BasicBlock.scala 132:19]
  wire  _GEN_62; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 716:29]
  assign _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 716:29]
  assign _T_6 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_6 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 727:32]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 75:58]
  assign predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 76:62]
  assign _T_14 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _T_15 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _T_16 = _T_14 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_17 = _T_15 | predicate_valid_R_1; // @[BasicBlock.scala 78:91]
  assign start = _T_16 & _T_17; // @[BasicBlock.scala 78:107]
  assign _T_22 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:52]
  assign _T_23 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_19 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_20 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_21 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_22 = start | _GEN_7; // @[BasicBlock.scala 112:19]
  assign _GEN_23 = start | _GEN_9; // @[BasicBlock.scala 112:19]
  assign _GEN_24 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_28 = {out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_29 = _T_28 == 4'hf; // @[HandShaking.scala 741:24]
  assign _T_32 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_33 = _T_32 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 726:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 715:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 715:21]
  assign io_Out_3_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 86:29]
  assign _GEN_54 = _T_23 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_55 = _GEN_54 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_56 = _GEN_55 & _T_29; // @[BasicBlock.scala 126:19]
  assign _GEN_57 = _GEN_56 & predicate; // @[BasicBlock.scala 126:19]
  assign _GEN_61 = predicate == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_62 = _GEN_56 & _GEN_61; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value = _RAND_9[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  state = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_23) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_29) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_23) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_29) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_23) begin
        if (_T_4) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_29) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_23) begin
        if (_T_5) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_29) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_23) begin
        out_valid_R_0 <= _GEN_19;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_23) begin
        out_valid_R_1 <= _GEN_20;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_23) begin
        out_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_4) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_23) begin
        out_valid_R_3 <= _GEN_22;
      end else begin
        if (_T_5) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_23) begin
        mask_valid_R_0 <= _GEN_23;
      end else begin
        if (_T_6) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_14) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_15) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_14) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_15) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_23) begin
        predicate_valid_R_0 <= _T_16;
      end else begin
        if (state) begin
          if (_T_29) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= _T_16;
          end
        end else begin
          predicate_valid_R_0 <= _T_16;
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_23) begin
        predicate_valid_R_1 <= _T_17;
      end else begin
        if (state) begin
          if (_T_29) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            predicate_valid_R_1 <= _T_17;
          end
        end else begin
          predicate_valid_R_1 <= _T_17;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_23) begin
        state <= _GEN_24;
      end else begin
        if (state) begin
          if (_T_29) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & _T_33) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body4: Output fired @ %d, Mask: %d\n",predicate_task,value,_T_22); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_62 & _T_33) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] bb_for_body4: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_4(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_6;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_7;
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_17; // @[BasicBlock.scala 309:81]
  wire  _T_18; // @[BasicBlock.scala 315:19]
  wire  _T_19; // @[BasicBlock.scala 315:19]
  wire  _GEN_6; // @[BasicBlock.scala 304:8]
  wire  _GEN_8; // @[BasicBlock.scala 304:8]
  wire  _GEN_26; // @[BasicBlock.scala 315:19]
  wire  _GEN_27; // @[BasicBlock.scala 315:19]
  wire  _GEN_29; // @[BasicBlock.scala 320:19]
  wire  _GEN_30; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_18 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_19 = _T_18 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_6 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_8 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_15 ? _GEN_6 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_26 = _T_15 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_27 = _GEN_26 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_29 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_17;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_8;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body7_preheader5: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body7_preheader5: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_5(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_6;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_7;
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_17; // @[BasicBlock.scala 309:81]
  wire  _T_18; // @[BasicBlock.scala 315:19]
  wire  _T_19; // @[BasicBlock.scala 315:19]
  wire  _GEN_6; // @[BasicBlock.scala 304:8]
  wire  _GEN_8; // @[BasicBlock.scala 304:8]
  wire  _GEN_26; // @[BasicBlock.scala 315:19]
  wire  _GEN_27; // @[BasicBlock.scala 315:19]
  wire  _GEN_29; // @[BasicBlock.scala 320:19]
  wire  _GEN_30; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_18 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_19 = _T_18 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_6 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_8 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_15 ? _GEN_6 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_26 = _T_15 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_27 = _GEN_26 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_29 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_17;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_8;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup6_loopexit6: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup6_loopexit6: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_6(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg [4:0] in_data_R_1_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_3;
  reg  in_data_R_1_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_4;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_5;
  reg  in_data_valid_R_1; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_6;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_7;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_8;
  reg  output_valid_R_1; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_9;
  reg  output_valid_R_2; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_10;
  reg  output_valid_R_3; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_11;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_12;
  reg  output_fire_R_1; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_13;
  reg  output_fire_R_2; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_14;
  reg  output_fire_R_3; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_15;
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[BasicBlock.scala 232:36]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 232:36]
  wire  _GEN_6; // @[BasicBlock.scala 232:36]
  wire [4:0] _T_11; // @[BasicBlock.scala 239:34]
  wire [4:0] _T_12; // @[BasicBlock.scala 239:34]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 240:15]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BasicBlock.scala 244:28]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BasicBlock.scala 244:28]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[BasicBlock.scala 244:28]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_1; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_2; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_3; // @[BasicBlock.scala 256:85]
  wire  predicate_val; // @[BasicBlock.scala 264:57]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_16;
  wire  _T_38; // @[Conditional.scala 37:30]
  wire  _T_39; // @[BasicBlock.scala 299:41]
  wire  _T_44; // @[BasicBlock.scala 309:81]
  wire  _T_45; // @[BasicBlock.scala 309:81]
  wire  _T_46; // @[BasicBlock.scala 309:81]
  wire  _T_47; // @[BasicBlock.scala 309:81]
  wire  _T_48; // @[BasicBlock.scala 315:19]
  wire  _T_49; // @[BasicBlock.scala 315:19]
  wire  _GEN_15; // @[BasicBlock.scala 304:8]
  wire  _GEN_16; // @[BasicBlock.scala 304:8]
  wire  _GEN_17; // @[BasicBlock.scala 304:8]
  wire  _GEN_18; // @[BasicBlock.scala 304:8]
  wire  _GEN_23; // @[BasicBlock.scala 304:8]
  wire  _T_53; // @[BasicBlock.scala 328:35]
  wire  _T_54; // @[BasicBlock.scala 328:35]
  wire  _T_55; // @[BasicBlock.scala 328:35]
  wire  _GEN_65; // @[BasicBlock.scala 315:19]
  wire  _GEN_66; // @[BasicBlock.scala 315:19]
  wire  _GEN_68; // @[BasicBlock.scala 320:19]
  wire  _GEN_69; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_8 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_8 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 232:36]
  assign _GEN_3 = _T_8 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign _T_10 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_10 ? io_predicateIn_1_bits_control : in_data_R_1_control; // @[BasicBlock.scala 232:36]
  assign _GEN_6 = _T_10 | in_data_valid_R_1; // @[BasicBlock.scala 232:36]
  assign _T_11 = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_12 = io_predicateIn_1_bits_taskID | in_data_R_1_taskID; // @[BasicBlock.scala 239:34]
  assign in_task_ID = _T_11 | _T_12; // @[BasicBlock.scala 240:15]
  assign _T_13 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_13 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign _T_14 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | output_fire_R_1; // @[BasicBlock.scala 244:28]
  assign _T_15 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_15 | output_fire_R_2; // @[BasicBlock.scala 244:28]
  assign _T_16 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | output_fire_R_3; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_13; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_1 = output_fire_R_1 | _T_14; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_2 = output_fire_R_2 | _T_15; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_3 = output_fire_R_3 | _T_16; // @[BasicBlock.scala 256:85]
  assign predicate_val = in_data_R_0_control | in_data_R_1_control; // @[BasicBlock.scala 264:57]
  assign _T_38 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_39 = _GEN_3 & _GEN_6; // @[BasicBlock.scala 299:41]
  assign _T_44 = _T_13 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_45 = _T_14 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_46 = _T_15 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_47 = _T_16 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_48 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_49 = _T_48 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_15 = _T_39 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_16 = _T_39 | output_valid_R_1; // @[BasicBlock.scala 304:8]
  assign _GEN_17 = _T_39 | output_valid_R_2; // @[BasicBlock.scala 304:8]
  assign _GEN_18 = _T_39 | output_valid_R_3; // @[BasicBlock.scala 304:8]
  assign _GEN_23 = _T_39 | state; // @[BasicBlock.scala 304:8]
  assign _T_53 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 328:35]
  assign _T_54 = _T_53 & out_fire_mask_2; // @[BasicBlock.scala 328:35]
  assign _T_55 = _T_54 & out_fire_mask_3; // @[BasicBlock.scala 328:35]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_predicateIn_1_ready = ~ in_data_valid_R_1; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_38 ? _GEN_15 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = _T_11 | _T_12; // @[BasicBlock.scala 282:22]
  assign io_Out_1_valid = _T_38 ? _GEN_16 : output_valid_R_1; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_1_bits_taskID = _T_11 | _T_12; // @[BasicBlock.scala 282:22]
  assign io_Out_1_bits_control = _GEN_1 | _GEN_4; // @[BasicBlock.scala 282:22]
  assign io_Out_2_valid = _T_38 ? _GEN_17 : output_valid_R_2; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_2_bits_taskID = _T_11 | _T_12; // @[BasicBlock.scala 282:22]
  assign io_Out_2_bits_control = _GEN_1 | _GEN_4; // @[BasicBlock.scala 282:22]
  assign io_Out_3_valid = _T_38 ? _GEN_18 : output_valid_R_3; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_3_bits_taskID = _T_11 | _T_12; // @[BasicBlock.scala 282:22]
  assign io_Out_3_bits_control = _GEN_1 | _GEN_4; // @[BasicBlock.scala 282:22]
  assign _GEN_65 = _T_38 & _T_39; // @[BasicBlock.scala 315:19]
  assign _GEN_66 = _GEN_65 & predicate_val; // @[BasicBlock.scala 315:19]
  assign _GEN_68 = predicate_val == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_69 = _GEN_65 & _GEN_68; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_R_1_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  state = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_38) begin
        if (_T_8) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_8) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_8) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_8) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_8) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_8) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_taskID <= 5'h0;
    end else begin
      if (_T_38) begin
        if (_T_10) begin
          in_data_R_1_taskID <= io_predicateIn_1_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_R_1_taskID <= 5'h0;
          end else begin
            if (_T_10) begin
              in_data_R_1_taskID <= io_predicateIn_1_bits_taskID;
            end
          end
        end else begin
          if (_T_10) begin
            in_data_R_1_taskID <= io_predicateIn_1_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_control <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_10) begin
          in_data_R_1_control <= io_predicateIn_1_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_R_1_control <= 1'h0;
          end else begin
            if (_T_10) begin
              in_data_R_1_control <= io_predicateIn_1_bits_control;
            end
          end
        end else begin
          if (_T_10) begin
            in_data_R_1_control <= io_predicateIn_1_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_38) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_38) begin
        in_data_valid_R_1 <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_6;
          end
        end else begin
          in_data_valid_R_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_39) begin
          output_valid_R_0 <= _T_44;
        end else begin
          if (_T_13) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_13) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_39) begin
          output_valid_R_1 <= _T_45;
        end else begin
          if (_T_14) begin
            output_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_14) begin
          output_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_39) begin
          output_valid_R_2 <= _T_46;
        end else begin
          if (_T_15) begin
            output_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_15) begin
          output_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_39) begin
          output_valid_R_3 <= _T_47;
        end else begin
          if (_T_16) begin
            output_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_16) begin
          output_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_38) begin
        output_fire_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_55) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_7;
          end
        end else begin
          output_fire_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else begin
      if (_T_38) begin
        output_fire_R_1 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_55) begin
            output_fire_R_1 <= 1'h0;
          end else begin
            output_fire_R_1 <= _GEN_9;
          end
        end else begin
          output_fire_R_1 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else begin
      if (_T_38) begin
        output_fire_R_2 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_55) begin
            output_fire_R_2 <= 1'h0;
          end else begin
            output_fire_R_2 <= _GEN_11;
          end
        end else begin
          output_fire_R_2 <= _GEN_11;
        end
      end
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else begin
      if (_T_38) begin
        output_fire_R_3 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_55) begin
            output_fire_R_3 <= 1'h0;
          end else begin
            output_fire_R_3 <= _GEN_13;
          end
        end else begin
          output_fire_R_3 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_38) begin
        state <= _GEN_23;
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & _T_49) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup67: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_49) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup67: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_1(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_2;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_3;
  reg  mask_valid_R_0; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_4;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 727:32]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_6;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_7;
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_8;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_9;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_10;
  reg  predicate_control_R_1; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_11;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_12;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_13;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_14;
  wire  predicate; // @[BasicBlock.scala 75:58]
  wire [4:0] predicate_task; // @[BasicBlock.scala 76:62]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _T_14; // @[BasicBlock.scala 78:91]
  wire  _T_15; // @[BasicBlock.scala 78:91]
  wire  start; // @[BasicBlock.scala 78:107]
  wire [1:0] _T_20; // @[BasicBlock.scala 102:52]
  wire  _T_21; // @[Conditional.scala 37:30]
  wire  _GEN_15; // @[BasicBlock.scala 112:19]
  wire  _GEN_16; // @[BasicBlock.scala 112:19]
  wire  _GEN_17; // @[BasicBlock.scala 112:19]
  wire  _GEN_18; // @[BasicBlock.scala 112:19]
  wire [1:0] _T_24; // @[HandShaking.scala 741:17]
  wire  _T_25; // @[HandShaking.scala 741:24]
  wire  _T_28; // @[BasicBlock.scala 126:19]
  wire  _T_29; // @[BasicBlock.scala 126:19]
  wire  _GEN_40; // @[BasicBlock.scala 126:19]
  wire  _GEN_41; // @[BasicBlock.scala 126:19]
  wire  _GEN_42; // @[BasicBlock.scala 126:19]
  wire  _GEN_43; // @[BasicBlock.scala 126:19]
  wire  _GEN_47; // @[BasicBlock.scala 132:19]
  wire  _GEN_48; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 727:32]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 75:58]
  assign predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 76:62]
  assign _T_12 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _T_13 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _T_14 = _T_12 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_15 = _T_13 | predicate_valid_R_1; // @[BasicBlock.scala 78:91]
  assign start = _T_14 & _T_15; // @[BasicBlock.scala 78:107]
  assign _T_20 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:52]
  assign _T_21 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_15 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_16 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_17 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_18 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_24 = {out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_25 = _T_24 == 2'h3; // @[HandShaking.scala 741:24]
  assign _T_28 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_29 = _T_28 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 726:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 86:29]
  assign _GEN_40 = _T_21 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_41 = _GEN_40 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_42 = _GEN_41 & _T_25; // @[BasicBlock.scala 126:19]
  assign _GEN_43 = _GEN_42 & predicate; // @[BasicBlock.scala 126:19]
  assign _GEN_47 = predicate == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_48 = _GEN_42 & _GEN_47; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_21) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_25) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_21) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_25) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_21) begin
        out_valid_R_0 <= _GEN_15;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_21) begin
        out_valid_R_1 <= _GEN_16;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_21) begin
        mask_valid_R_0 <= _GEN_17;
      end else begin
        if (_T_4) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_12) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_13) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_13) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_13) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_21) begin
        predicate_valid_R_0 <= _T_14;
      end else begin
        if (state) begin
          if (_T_25) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= _T_14;
          end
        end else begin
          predicate_valid_R_0 <= _T_14;
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_21) begin
        predicate_valid_R_1 <= _T_15;
      end else begin
        if (state) begin
          if (_T_25) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            predicate_valid_R_1 <= _T_15;
          end
        end else begin
          predicate_valid_R_1 <= _T_15;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_21) begin
        state <= _GEN_18;
      end else begin
        if (state) begin
          if (_T_25) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_43 & _T_29) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body78: Output fired @ %d, Mask: %d\n",predicate_task,value,_T_20); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_48 & _T_29) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] bb_for_body78: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_7(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_valid_R_1; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_6;
  reg  output_valid_R_2; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_7;
  reg  output_valid_R_3; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_8;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_9;
  reg  output_fire_R_1; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_10;
  reg  output_fire_R_2; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_11;
  reg  output_fire_R_3; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_12;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BasicBlock.scala 244:28]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[BasicBlock.scala 244:28]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_10; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_1; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_2; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_3; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_13;
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _T_29; // @[BasicBlock.scala 309:81]
  wire  _T_30; // @[BasicBlock.scala 309:81]
  wire  _T_31; // @[BasicBlock.scala 309:81]
  wire  _T_32; // @[BasicBlock.scala 309:81]
  wire  _T_33; // @[BasicBlock.scala 315:19]
  wire  _T_34; // @[BasicBlock.scala 315:19]
  wire  _GEN_12; // @[BasicBlock.scala 304:8]
  wire  _GEN_13; // @[BasicBlock.scala 304:8]
  wire  _GEN_14; // @[BasicBlock.scala 304:8]
  wire  _GEN_15; // @[BasicBlock.scala 304:8]
  wire  _GEN_20; // @[BasicBlock.scala 304:8]
  wire  _T_38; // @[BasicBlock.scala 328:35]
  wire  _T_39; // @[BasicBlock.scala 328:35]
  wire  _T_40; // @[BasicBlock.scala 328:35]
  wire  _GEN_53; // @[BasicBlock.scala 315:19]
  wire  _GEN_54; // @[BasicBlock.scala 315:19]
  wire  _GEN_56; // @[BasicBlock.scala 320:19]
  wire  _GEN_57; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 244:28]
  assign _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 244:28]
  assign _T_11 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_10 = _T_11 | output_fire_R_3; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_3 = output_fire_R_3 | _T_11; // @[BasicBlock.scala 256:85]
  assign _T_24 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_29 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_30 = _T_9 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_31 = _T_10 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_32 = _T_11 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_33 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_34 = _T_33 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_12 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_13 = _GEN_3 | output_valid_R_1; // @[BasicBlock.scala 304:8]
  assign _GEN_14 = _GEN_3 | output_valid_R_2; // @[BasicBlock.scala 304:8]
  assign _GEN_15 = _GEN_3 | output_valid_R_3; // @[BasicBlock.scala 304:8]
  assign _GEN_20 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign _T_38 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 328:35]
  assign _T_39 = _T_38 & out_fire_mask_2; // @[BasicBlock.scala 328:35]
  assign _T_40 = _T_39 & out_fire_mask_3; // @[BasicBlock.scala 328:35]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_24 ? _GEN_12 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_1_valid = _T_24 ? _GEN_13 : output_valid_R_1; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_1_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_2_valid = _T_24 ? _GEN_14 : output_valid_R_2; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_2_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_3_valid = _T_24 ? _GEN_15 : output_valid_R_3; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_3_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_3_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_53 = _T_24 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_54 = _GEN_53 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_56 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_57 = _GEN_53 & _GEN_56; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  state = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_24) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_40) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_40) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_40) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_29;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_GEN_3) begin
          output_valid_R_1 <= _T_30;
        end else begin
          if (_T_9) begin
            output_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_9) begin
          output_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_GEN_3) begin
          output_valid_R_2 <= _T_31;
        end else begin
          if (_T_10) begin
            output_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_10) begin
          output_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_GEN_3) begin
          output_valid_R_3 <= _T_32;
        end else begin
          if (_T_11) begin
            output_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_11) begin
          output_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (_T_40) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        output_fire_R_1 <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_40) begin
            output_fire_R_1 <= 1'h0;
          end else begin
            output_fire_R_1 <= _GEN_6;
          end
        end else begin
          output_fire_R_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        output_fire_R_2 <= _GEN_8;
      end else begin
        if (state) begin
          if (_T_40) begin
            output_fire_R_2 <= 1'h0;
          end else begin
            output_fire_R_2 <= _GEN_8;
          end
        end else begin
          output_fire_R_2 <= _GEN_8;
        end
      end
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        output_fire_R_3 <= _GEN_10;
      end else begin
        if (state) begin
          if (_T_40) begin
            output_fire_R_3 <= 1'h0;
          end else begin
            output_fire_R_3 <= _GEN_10;
          end
        end else begin
          output_fire_R_3 <= _GEN_10;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_24) begin
        state <= _GEN_20;
      end else begin
        if (state) begin
          if (_T_40) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_54 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body15_lr_ph9: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body15_lr_ph9: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_8(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_6;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_7;
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_17; // @[BasicBlock.scala 309:81]
  wire  _T_18; // @[BasicBlock.scala 315:19]
  wire  _T_19; // @[BasicBlock.scala 315:19]
  wire  _GEN_6; // @[BasicBlock.scala 304:8]
  wire  _GEN_8; // @[BasicBlock.scala 304:8]
  wire  _GEN_26; // @[BasicBlock.scala 315:19]
  wire  _GEN_27; // @[BasicBlock.scala 315:19]
  wire  _GEN_29; // @[BasicBlock.scala 320:19]
  wire  _GEN_30; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_18 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_19 = _T_18 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_6 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_8 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_15 ? _GEN_6 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_26 = _T_15 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_27 = _GEN_26 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_29 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_17;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_8;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup14_loopexit10: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup14_loopexit10: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_9(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg [4:0] in_data_R_1_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_3;
  reg  in_data_R_1_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_4;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_5;
  reg  in_data_valid_R_1; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_6;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_7;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_8;
  reg  output_valid_R_1; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_9;
  reg  output_valid_R_2; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_10;
  reg  output_valid_R_3; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_11;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_12;
  reg  output_fire_R_1; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_13;
  reg  output_fire_R_2; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_14;
  reg  output_fire_R_3; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_15;
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[BasicBlock.scala 232:36]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 232:36]
  wire  _GEN_6; // @[BasicBlock.scala 232:36]
  wire [4:0] _T_11; // @[BasicBlock.scala 239:34]
  wire [4:0] _T_12; // @[BasicBlock.scala 239:34]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 240:15]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BasicBlock.scala 244:28]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BasicBlock.scala 244:28]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[BasicBlock.scala 244:28]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_1; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_2; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_3; // @[BasicBlock.scala 256:85]
  wire  predicate_val; // @[BasicBlock.scala 264:57]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_16;
  wire  _T_38; // @[Conditional.scala 37:30]
  wire  _T_39; // @[BasicBlock.scala 299:41]
  wire  _T_44; // @[BasicBlock.scala 309:81]
  wire  _T_45; // @[BasicBlock.scala 309:81]
  wire  _T_46; // @[BasicBlock.scala 309:81]
  wire  _T_47; // @[BasicBlock.scala 309:81]
  wire  _T_48; // @[BasicBlock.scala 315:19]
  wire  _T_49; // @[BasicBlock.scala 315:19]
  wire  _GEN_15; // @[BasicBlock.scala 304:8]
  wire  _GEN_16; // @[BasicBlock.scala 304:8]
  wire  _GEN_17; // @[BasicBlock.scala 304:8]
  wire  _GEN_18; // @[BasicBlock.scala 304:8]
  wire  _GEN_23; // @[BasicBlock.scala 304:8]
  wire  _T_53; // @[BasicBlock.scala 328:35]
  wire  _T_54; // @[BasicBlock.scala 328:35]
  wire  _T_55; // @[BasicBlock.scala 328:35]
  wire  _GEN_65; // @[BasicBlock.scala 315:19]
  wire  _GEN_66; // @[BasicBlock.scala 315:19]
  wire  _GEN_68; // @[BasicBlock.scala 320:19]
  wire  _GEN_69; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_8 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_8 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 232:36]
  assign _GEN_3 = _T_8 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign _T_10 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_10 ? io_predicateIn_1_bits_control : in_data_R_1_control; // @[BasicBlock.scala 232:36]
  assign _GEN_6 = _T_10 | in_data_valid_R_1; // @[BasicBlock.scala 232:36]
  assign _T_11 = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_12 = io_predicateIn_1_bits_taskID | in_data_R_1_taskID; // @[BasicBlock.scala 239:34]
  assign in_task_ID = _T_11 | _T_12; // @[BasicBlock.scala 240:15]
  assign _T_13 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_13 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign _T_14 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | output_fire_R_1; // @[BasicBlock.scala 244:28]
  assign _T_15 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_15 | output_fire_R_2; // @[BasicBlock.scala 244:28]
  assign _T_16 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | output_fire_R_3; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_13; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_1 = output_fire_R_1 | _T_14; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_2 = output_fire_R_2 | _T_15; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_3 = output_fire_R_3 | _T_16; // @[BasicBlock.scala 256:85]
  assign predicate_val = in_data_R_0_control | in_data_R_1_control; // @[BasicBlock.scala 264:57]
  assign _T_38 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_39 = _GEN_3 & _GEN_6; // @[BasicBlock.scala 299:41]
  assign _T_44 = _T_13 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_45 = _T_14 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_46 = _T_15 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_47 = _T_16 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_48 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_49 = _T_48 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_15 = _T_39 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_16 = _T_39 | output_valid_R_1; // @[BasicBlock.scala 304:8]
  assign _GEN_17 = _T_39 | output_valid_R_2; // @[BasicBlock.scala 304:8]
  assign _GEN_18 = _T_39 | output_valid_R_3; // @[BasicBlock.scala 304:8]
  assign _GEN_23 = _T_39 | state; // @[BasicBlock.scala 304:8]
  assign _T_53 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 328:35]
  assign _T_54 = _T_53 & out_fire_mask_2; // @[BasicBlock.scala 328:35]
  assign _T_55 = _T_54 & out_fire_mask_3; // @[BasicBlock.scala 328:35]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_predicateIn_1_ready = ~ in_data_valid_R_1; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_38 ? _GEN_15 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = _T_11 | _T_12; // @[BasicBlock.scala 282:22]
  assign io_Out_1_valid = _T_38 ? _GEN_16 : output_valid_R_1; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_1_bits_taskID = _T_11 | _T_12; // @[BasicBlock.scala 282:22]
  assign io_Out_1_bits_control = _GEN_1 | _GEN_4; // @[BasicBlock.scala 282:22]
  assign io_Out_2_valid = _T_38 ? _GEN_17 : output_valid_R_2; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_2_bits_taskID = _T_11 | _T_12; // @[BasicBlock.scala 282:22]
  assign io_Out_2_bits_control = _GEN_1 | _GEN_4; // @[BasicBlock.scala 282:22]
  assign io_Out_3_valid = _T_38 ? _GEN_18 : output_valid_R_3; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_3_bits_taskID = _T_11 | _T_12; // @[BasicBlock.scala 282:22]
  assign io_Out_3_bits_control = _GEN_1 | _GEN_4; // @[BasicBlock.scala 282:22]
  assign _GEN_65 = _T_38 & _T_39; // @[BasicBlock.scala 315:19]
  assign _GEN_66 = _GEN_65 & predicate_val; // @[BasicBlock.scala 315:19]
  assign _GEN_68 = predicate_val == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_69 = _GEN_65 & _GEN_68; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_R_1_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  state = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_38) begin
        if (_T_8) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_8) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_8) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_8) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_8) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_8) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_taskID <= 5'h0;
    end else begin
      if (_T_38) begin
        if (_T_10) begin
          in_data_R_1_taskID <= io_predicateIn_1_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_R_1_taskID <= 5'h0;
          end else begin
            if (_T_10) begin
              in_data_R_1_taskID <= io_predicateIn_1_bits_taskID;
            end
          end
        end else begin
          if (_T_10) begin
            in_data_R_1_taskID <= io_predicateIn_1_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_control <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_10) begin
          in_data_R_1_control <= io_predicateIn_1_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_R_1_control <= 1'h0;
          end else begin
            if (_T_10) begin
              in_data_R_1_control <= io_predicateIn_1_bits_control;
            end
          end
        end else begin
          if (_T_10) begin
            in_data_R_1_control <= io_predicateIn_1_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_38) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_38) begin
        in_data_valid_R_1 <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_55) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_6;
          end
        end else begin
          in_data_valid_R_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_39) begin
          output_valid_R_0 <= _T_44;
        end else begin
          if (_T_13) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_13) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_39) begin
          output_valid_R_1 <= _T_45;
        end else begin
          if (_T_14) begin
            output_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_14) begin
          output_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_39) begin
          output_valid_R_2 <= _T_46;
        end else begin
          if (_T_15) begin
            output_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_15) begin
          output_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else begin
      if (_T_38) begin
        if (_T_39) begin
          output_valid_R_3 <= _T_47;
        end else begin
          if (_T_16) begin
            output_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_16) begin
          output_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_38) begin
        output_fire_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_55) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_7;
          end
        end else begin
          output_fire_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else begin
      if (_T_38) begin
        output_fire_R_1 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_55) begin
            output_fire_R_1 <= 1'h0;
          end else begin
            output_fire_R_1 <= _GEN_9;
          end
        end else begin
          output_fire_R_1 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else begin
      if (_T_38) begin
        output_fire_R_2 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_55) begin
            output_fire_R_2 <= 1'h0;
          end else begin
            output_fire_R_2 <= _GEN_11;
          end
        end else begin
          output_fire_R_2 <= _GEN_11;
        end
      end
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else begin
      if (_T_38) begin
        output_fire_R_3 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_55) begin
            output_fire_R_3 <= 1'h0;
          end else begin
            output_fire_R_3 <= _GEN_13;
          end
        end else begin
          output_fire_R_3 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_38) begin
        state <= _GEN_23;
      end else begin
        if (state) begin
          if (_T_55) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & _T_49) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup1411: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_49) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup1411: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_2(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output       io_Out_0_bits_control,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output [4:0] io_Out_5_bits_taskID,
  output       io_Out_5_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_4;
  reg  out_ready_R_5; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_5;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_6;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_7;
  reg  out_valid_R_2; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_8;
  reg  out_valid_R_3; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_9;
  reg  out_valid_R_4; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_10;
  reg  out_valid_R_5; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_11;
  reg  mask_valid_R_0; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_12;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 716:29]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[HandShaking.scala 716:29]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[HandShaking.scala 716:29]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[HandShaking.scala 716:29]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[HandShaking.scala 727:32]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_13;
  wire [14:0] _T_11; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_14;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_15;
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_16;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_17;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_18;
  reg  predicate_control_R_1; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_19;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_20;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_21;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_22;
  wire  predicate; // @[BasicBlock.scala 75:58]
  wire [4:0] predicate_task; // @[BasicBlock.scala 76:62]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _T_17; // @[Decoupled.scala 40:37]
  wire  _T_18; // @[BasicBlock.scala 78:91]
  wire  _T_19; // @[BasicBlock.scala 78:91]
  wire  start; // @[BasicBlock.scala 78:107]
  wire [1:0] _T_24; // @[BasicBlock.scala 102:52]
  wire  _T_25; // @[Conditional.scala 37:30]
  wire  _GEN_23; // @[BasicBlock.scala 112:19]
  wire  _GEN_24; // @[BasicBlock.scala 112:19]
  wire  _GEN_25; // @[BasicBlock.scala 112:19]
  wire  _GEN_26; // @[BasicBlock.scala 112:19]
  wire  _GEN_27; // @[BasicBlock.scala 112:19]
  wire  _GEN_28; // @[BasicBlock.scala 112:19]
  wire  _GEN_29; // @[BasicBlock.scala 112:19]
  wire  _GEN_30; // @[BasicBlock.scala 112:19]
  wire [5:0] _T_32; // @[HandShaking.scala 741:17]
  wire  _T_33; // @[HandShaking.scala 741:24]
  wire  _T_36; // @[BasicBlock.scala 126:19]
  wire  _T_37; // @[BasicBlock.scala 126:19]
  wire  _GEN_68; // @[BasicBlock.scala 126:19]
  wire  _GEN_69; // @[BasicBlock.scala 126:19]
  wire  _GEN_70; // @[BasicBlock.scala 126:19]
  wire  _GEN_71; // @[BasicBlock.scala 126:19]
  wire  _GEN_75; // @[BasicBlock.scala 132:19]
  wire  _GEN_76; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 716:29]
  assign _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 716:29]
  assign _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 716:29]
  assign _T_7 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_7 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 716:29]
  assign _T_8 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_8 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 727:32]
  assign _T_11 = value + 15'h1; // @[Counter.scala 38:22]
  assign predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 75:58]
  assign predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 76:62]
  assign _T_16 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _T_17 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _T_18 = _T_16 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_19 = _T_17 | predicate_valid_R_1; // @[BasicBlock.scala 78:91]
  assign start = _T_18 & _T_19; // @[BasicBlock.scala 78:107]
  assign _T_24 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:52]
  assign _T_25 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_23 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_24 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_25 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_26 = start | _GEN_7; // @[BasicBlock.scala 112:19]
  assign _GEN_27 = start | _GEN_9; // @[BasicBlock.scala 112:19]
  assign _GEN_28 = start | _GEN_11; // @[BasicBlock.scala 112:19]
  assign _GEN_29 = start | _GEN_13; // @[BasicBlock.scala 112:19]
  assign _GEN_30 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_32 = {out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_33 = _T_32 == 6'h3f; // @[HandShaking.scala 741:24]
  assign _T_36 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_37 = _T_36 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 726:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 715:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 715:21]
  assign io_Out_3_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 715:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 715:21]
  assign io_Out_5_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_5_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 86:29]
  assign _GEN_68 = _T_25 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_69 = _GEN_68 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_70 = _GEN_69 & _T_33; // @[BasicBlock.scala 126:19]
  assign _GEN_71 = _GEN_70 & predicate; // @[BasicBlock.scala 126:19]
  assign _GEN_75 = predicate == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_76 = _GEN_70 & _GEN_75; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  value = _RAND_13[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  state = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_25) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_33) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_25) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_33) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_25) begin
        if (_T_4) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_33) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_25) begin
        if (_T_5) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_33) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_25) begin
        if (_T_6) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_33) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_6) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_6) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_25) begin
        if (_T_7) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_33) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_7) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_7) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_25) begin
        out_valid_R_0 <= _GEN_23;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_25) begin
        out_valid_R_1 <= _GEN_24;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_25) begin
        out_valid_R_2 <= _GEN_25;
      end else begin
        if (_T_4) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_25) begin
        out_valid_R_3 <= _GEN_26;
      end else begin
        if (_T_5) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_25) begin
        out_valid_R_4 <= _GEN_27;
      end else begin
        if (_T_6) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_25) begin
        out_valid_R_5 <= _GEN_28;
      end else begin
        if (_T_7) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_25) begin
        mask_valid_R_0 <= _GEN_29;
      end else begin
        if (_T_8) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_11;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_16) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_16) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_17) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_17) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_25) begin
        predicate_valid_R_0 <= _T_18;
      end else begin
        if (state) begin
          if (_T_33) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= _T_18;
          end
        end else begin
          predicate_valid_R_0 <= _T_18;
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_25) begin
        predicate_valid_R_1 <= _T_19;
      end else begin
        if (state) begin
          if (_T_33) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            predicate_valid_R_1 <= _T_19;
          end
        end else begin
          predicate_valid_R_1 <= _T_19;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_25) begin
        state <= _GEN_30;
      end else begin
        if (state) begin
          if (_T_33) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & _T_37) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body1512: Output fired @ %d, Mask: %d\n",predicate_task,value,_T_24); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_76 & _T_37) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] bb_for_body1512: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_10(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_valid_R_1; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_6;
  reg  output_valid_R_2; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_7;
  reg  output_valid_R_3; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_8;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_9;
  reg  output_fire_R_1; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_10;
  reg  output_fire_R_2; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_11;
  reg  output_fire_R_3; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_12;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BasicBlock.scala 244:28]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[BasicBlock.scala 244:28]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_10; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_1; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_2; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_3; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_13;
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _T_29; // @[BasicBlock.scala 309:81]
  wire  _T_30; // @[BasicBlock.scala 309:81]
  wire  _T_31; // @[BasicBlock.scala 309:81]
  wire  _T_32; // @[BasicBlock.scala 309:81]
  wire  _T_33; // @[BasicBlock.scala 315:19]
  wire  _T_34; // @[BasicBlock.scala 315:19]
  wire  _GEN_12; // @[BasicBlock.scala 304:8]
  wire  _GEN_13; // @[BasicBlock.scala 304:8]
  wire  _GEN_14; // @[BasicBlock.scala 304:8]
  wire  _GEN_15; // @[BasicBlock.scala 304:8]
  wire  _GEN_20; // @[BasicBlock.scala 304:8]
  wire  _T_38; // @[BasicBlock.scala 328:35]
  wire  _T_39; // @[BasicBlock.scala 328:35]
  wire  _T_40; // @[BasicBlock.scala 328:35]
  wire  _GEN_53; // @[BasicBlock.scala 315:19]
  wire  _GEN_54; // @[BasicBlock.scala 315:19]
  wire  _GEN_56; // @[BasicBlock.scala 320:19]
  wire  _GEN_57; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 244:28]
  assign _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 244:28]
  assign _T_11 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_10 = _T_11 | output_fire_R_3; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_3 = output_fire_R_3 | _T_11; // @[BasicBlock.scala 256:85]
  assign _T_24 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_29 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_30 = _T_9 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_31 = _T_10 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_32 = _T_11 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_33 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_34 = _T_33 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_12 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_13 = _GEN_3 | output_valid_R_1; // @[BasicBlock.scala 304:8]
  assign _GEN_14 = _GEN_3 | output_valid_R_2; // @[BasicBlock.scala 304:8]
  assign _GEN_15 = _GEN_3 | output_valid_R_3; // @[BasicBlock.scala 304:8]
  assign _GEN_20 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign _T_38 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 328:35]
  assign _T_39 = _T_38 & out_fire_mask_2; // @[BasicBlock.scala 328:35]
  assign _T_40 = _T_39 & out_fire_mask_3; // @[BasicBlock.scala 328:35]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_24 ? _GEN_12 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_1_valid = _T_24 ? _GEN_13 : output_valid_R_1; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_1_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_2_valid = _T_24 ? _GEN_14 : output_valid_R_2; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_2_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_3_valid = _T_24 ? _GEN_15 : output_valid_R_3; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_3_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_3_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_53 = _T_24 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_54 = _GEN_53 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_56 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_57 = _GEN_53 & _GEN_56; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  state = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_24) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_40) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_40) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_40) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_29;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_GEN_3) begin
          output_valid_R_1 <= _T_30;
        end else begin
          if (_T_9) begin
            output_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_9) begin
          output_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_GEN_3) begin
          output_valid_R_2 <= _T_31;
        end else begin
          if (_T_10) begin
            output_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_10) begin
          output_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_GEN_3) begin
          output_valid_R_3 <= _T_32;
        end else begin
          if (_T_11) begin
            output_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_11) begin
          output_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (_T_40) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        output_fire_R_1 <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_40) begin
            output_fire_R_1 <= 1'h0;
          end else begin
            output_fire_R_1 <= _GEN_6;
          end
        end else begin
          output_fire_R_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        output_fire_R_2 <= _GEN_8;
      end else begin
        if (state) begin
          if (_T_40) begin
            output_fire_R_2 <= 1'h0;
          end else begin
            output_fire_R_2 <= _GEN_8;
          end
        end else begin
          output_fire_R_2 <= _GEN_8;
        end
      end
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        output_fire_R_3 <= _GEN_10;
      end else begin
        if (state) begin
          if (_T_40) begin
            output_fire_R_3 <= 1'h0;
          end else begin
            output_fire_R_3 <= _GEN_10;
          end
        end else begin
          output_fire_R_3 <= _GEN_10;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_24) begin
        state <= _GEN_20;
      end else begin
        if (state) begin
          if (_T_40) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_54 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup2013: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_57 & _T_34) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup2013: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_3(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output       io_Out_1_bits_control,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_6;
  reg  out_valid_R_2; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_7;
  reg  out_valid_R_3; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_8;
  reg  out_valid_R_4; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_9;
  reg  mask_valid_R_0; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_10;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 716:29]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[HandShaking.scala 716:29]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[HandShaking.scala 716:29]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[HandShaking.scala 727:32]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_11;
  wire [14:0] _T_10; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_12;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_13;
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_14;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_15;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_16;
  reg  predicate_control_R_1; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_17;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_18;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_19;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_20;
  wire  predicate; // @[BasicBlock.scala 75:58]
  wire [4:0] predicate_task; // @[BasicBlock.scala 76:62]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _T_17; // @[BasicBlock.scala 78:91]
  wire  _T_18; // @[BasicBlock.scala 78:91]
  wire  start; // @[BasicBlock.scala 78:107]
  wire [1:0] _T_23; // @[BasicBlock.scala 102:52]
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _GEN_21; // @[BasicBlock.scala 112:19]
  wire  _GEN_22; // @[BasicBlock.scala 112:19]
  wire  _GEN_23; // @[BasicBlock.scala 112:19]
  wire  _GEN_24; // @[BasicBlock.scala 112:19]
  wire  _GEN_25; // @[BasicBlock.scala 112:19]
  wire  _GEN_26; // @[BasicBlock.scala 112:19]
  wire  _GEN_27; // @[BasicBlock.scala 112:19]
  wire [4:0] _T_30; // @[HandShaking.scala 741:17]
  wire  _T_31; // @[HandShaking.scala 741:24]
  wire  _T_34; // @[BasicBlock.scala 126:19]
  wire  _T_35; // @[BasicBlock.scala 126:19]
  wire  _GEN_61; // @[BasicBlock.scala 126:19]
  wire  _GEN_62; // @[BasicBlock.scala 126:19]
  wire  _GEN_63; // @[BasicBlock.scala 126:19]
  wire  _GEN_64; // @[BasicBlock.scala 126:19]
  wire  _GEN_68; // @[BasicBlock.scala 132:19]
  wire  _GEN_69; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 716:29]
  assign _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 716:29]
  assign _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 716:29]
  assign _T_7 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_7 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 727:32]
  assign _T_10 = value + 15'h1; // @[Counter.scala 38:22]
  assign predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 75:58]
  assign predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 76:62]
  assign _T_15 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _T_16 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _T_17 = _T_15 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_18 = _T_16 | predicate_valid_R_1; // @[BasicBlock.scala 78:91]
  assign start = _T_17 & _T_18; // @[BasicBlock.scala 78:107]
  assign _T_23 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:52]
  assign _T_24 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_21 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_22 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_23 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_24 = start | _GEN_7; // @[BasicBlock.scala 112:19]
  assign _GEN_25 = start | _GEN_9; // @[BasicBlock.scala 112:19]
  assign _GEN_26 = start | _GEN_11; // @[BasicBlock.scala 112:19]
  assign _GEN_27 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_30 = {out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_31 = _T_30 == 5'h1f; // @[HandShaking.scala 741:24]
  assign _T_34 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_35 = _T_34 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 726:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 715:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 715:21]
  assign io_Out_3_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 715:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 86:29]
  assign _GEN_61 = _T_24 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_62 = _GEN_61 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_63 = _GEN_62 & _T_31; // @[BasicBlock.scala 126:19]
  assign _GEN_64 = _GEN_63 & predicate; // @[BasicBlock.scala 126:19]
  assign _GEN_68 = predicate == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_69 = _GEN_63 & _GEN_68; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  value = _RAND_11[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_12[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  state = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_31) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_31) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_4) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_31) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_5) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_31) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_6) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_31) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_6) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_6) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_0 <= _GEN_21;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_1 <= _GEN_22;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_2 <= _GEN_23;
      end else begin
        if (_T_4) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_3 <= _GEN_24;
      end else begin
        if (_T_5) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_4 <= _GEN_25;
      end else begin
        if (_T_6) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        mask_valid_R_0 <= _GEN_26;
      end else begin
        if (_T_7) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_10;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_15) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_16) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_16) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_16) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        predicate_valid_R_0 <= _T_17;
      end else begin
        if (state) begin
          if (_T_31) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= _T_17;
          end
        end else begin
          predicate_valid_R_0 <= _T_17;
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        predicate_valid_R_1 <= _T_18;
      end else begin
        if (state) begin
          if (_T_31) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            predicate_valid_R_1 <= _T_18;
          end
        end else begin
          predicate_valid_R_1 <= _T_18;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_24) begin
        state <= _GEN_27;
      end else begin
        if (state) begin
          if (_T_31) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_64 & _T_35) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body2114: Output fired @ %d, Mask: %d\n",predicate_task,value,_T_23); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_35) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] bb_for_body2114: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_4(
  input        clock,
  input        reset,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output [4:0] io_Out_5_bits_taskID,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output [4:0] io_Out_6_bits_taskID,
  output       io_Out_6_bits_control,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output [4:0] io_Out_7_bits_taskID,
  output       io_Out_7_bits_control,
  input        io_Out_8_ready,
  output       io_Out_8_valid,
  output [4:0] io_Out_8_bits_taskID,
  output       io_Out_8_bits_control,
  input        io_Out_9_ready,
  output       io_Out_9_valid,
  output [4:0] io_Out_9_bits_taskID,
  output       io_Out_9_bits_control,
  input        io_Out_10_ready,
  output       io_Out_10_valid,
  output [4:0] io_Out_10_bits_taskID,
  output       io_Out_10_bits_control,
  input        io_Out_11_ready,
  output       io_Out_11_valid,
  output [4:0] io_Out_11_bits_taskID,
  output       io_Out_11_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_4;
  reg  out_ready_R_5; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_5;
  reg  out_ready_R_6; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_6;
  reg  out_ready_R_7; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_7;
  reg  out_ready_R_8; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_8;
  reg  out_ready_R_9; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_9;
  reg  out_ready_R_10; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_10;
  reg  out_ready_R_11; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_11;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_12;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_13;
  reg  out_valid_R_2; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_14;
  reg  out_valid_R_3; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_15;
  reg  out_valid_R_4; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_16;
  reg  out_valid_R_5; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_17;
  reg  out_valid_R_6; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_18;
  reg  out_valid_R_7; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_19;
  reg  out_valid_R_8; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_20;
  reg  out_valid_R_9; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_21;
  reg  out_valid_R_10; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_22;
  reg  out_valid_R_11; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_23;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 716:29]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[HandShaking.scala 716:29]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[HandShaking.scala 716:29]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[HandShaking.scala 716:29]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[HandShaking.scala 716:29]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[HandShaking.scala 716:29]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[HandShaking.scala 716:29]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[HandShaking.scala 716:29]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[HandShaking.scala 716:29]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_23; // @[HandShaking.scala 716:29]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_24;
  wire [14:0] _T_17; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_25;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_26;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_27;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_28;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_29;
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  start; // @[BasicBlock.scala 78:91]
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _GEN_31; // @[BasicBlock.scala 112:19]
  wire  _GEN_32; // @[BasicBlock.scala 112:19]
  wire  _GEN_33; // @[BasicBlock.scala 112:19]
  wire  _GEN_34; // @[BasicBlock.scala 112:19]
  wire  _GEN_35; // @[BasicBlock.scala 112:19]
  wire  _GEN_36; // @[BasicBlock.scala 112:19]
  wire  _GEN_37; // @[BasicBlock.scala 112:19]
  wire  _GEN_38; // @[BasicBlock.scala 112:19]
  wire  _GEN_39; // @[BasicBlock.scala 112:19]
  wire  _GEN_40; // @[BasicBlock.scala 112:19]
  wire  _GEN_41; // @[BasicBlock.scala 112:19]
  wire  _GEN_42; // @[BasicBlock.scala 112:19]
  wire  _GEN_44; // @[BasicBlock.scala 112:19]
  wire [5:0] _T_31; // @[HandShaking.scala 741:17]
  wire [11:0] _T_37; // @[HandShaking.scala 741:17]
  wire  _T_38; // @[HandShaking.scala 741:24]
  wire  _T_40; // @[BasicBlock.scala 126:19]
  wire  _T_41; // @[BasicBlock.scala 126:19]
  wire  _GEN_103; // @[BasicBlock.scala 126:19]
  wire  _GEN_104; // @[BasicBlock.scala 126:19]
  wire  _GEN_105; // @[BasicBlock.scala 126:19]
  wire  _GEN_106; // @[BasicBlock.scala 126:19]
  wire  _GEN_110; // @[BasicBlock.scala 132:19]
  wire  _GEN_111; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 716:29]
  assign _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 716:29]
  assign _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 716:29]
  assign _T_7 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_7 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 716:29]
  assign _T_8 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_8 ? 1'h0 : out_valid_R_6; // @[HandShaking.scala 716:29]
  assign _T_9 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_9 ? 1'h0 : out_valid_R_7; // @[HandShaking.scala 716:29]
  assign _T_10 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_10 ? 1'h0 : out_valid_R_8; // @[HandShaking.scala 716:29]
  assign _T_11 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_11 ? 1'h0 : out_valid_R_9; // @[HandShaking.scala 716:29]
  assign _T_12 = io_Out_10_ready & io_Out_10_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_12 ? 1'h0 : out_valid_R_10; // @[HandShaking.scala 716:29]
  assign _T_13 = io_Out_11_ready & io_Out_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_23 = _T_13 ? 1'h0 : out_valid_R_11; // @[HandShaking.scala 716:29]
  assign _T_17 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_21 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign start = _T_21 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_24 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_31 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_32 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_33 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_34 = start | _GEN_7; // @[BasicBlock.scala 112:19]
  assign _GEN_35 = start | _GEN_9; // @[BasicBlock.scala 112:19]
  assign _GEN_36 = start | _GEN_11; // @[BasicBlock.scala 112:19]
  assign _GEN_37 = start | _GEN_13; // @[BasicBlock.scala 112:19]
  assign _GEN_38 = start | _GEN_15; // @[BasicBlock.scala 112:19]
  assign _GEN_39 = start | _GEN_17; // @[BasicBlock.scala 112:19]
  assign _GEN_40 = start | _GEN_19; // @[BasicBlock.scala 112:19]
  assign _GEN_41 = start | _GEN_21; // @[BasicBlock.scala 112:19]
  assign _GEN_42 = start | _GEN_23; // @[BasicBlock.scala 112:19]
  assign _GEN_44 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_31 = {out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_37 = {out_ready_R_11,out_ready_R_10,out_ready_R_9,out_ready_R_8,out_ready_R_7,out_ready_R_6,_T_31}; // @[HandShaking.scala 741:17]
  assign _T_38 = _T_37 == 12'hfff; // @[HandShaking.scala 741:24]
  assign _T_40 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_41 = _T_40 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 715:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 715:21]
  assign io_Out_3_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 715:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_4_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 715:21]
  assign io_Out_5_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 715:21]
  assign io_Out_6_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_6_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 715:21]
  assign io_Out_7_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_7_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_8_valid = out_valid_R_8; // @[HandShaking.scala 715:21]
  assign io_Out_8_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_8_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_9_valid = out_valid_R_9; // @[HandShaking.scala 715:21]
  assign io_Out_9_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_9_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_10_valid = out_valid_R_10; // @[HandShaking.scala 715:21]
  assign io_Out_10_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_10_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_11_valid = out_valid_R_11; // @[HandShaking.scala 715:21]
  assign io_Out_11_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_11_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign _GEN_103 = _T_24 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_104 = _GEN_103 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_105 = _GEN_104 & _T_38; // @[BasicBlock.scala 126:19]
  assign _GEN_106 = _GEN_105 & predicate_in_R_0_control; // @[BasicBlock.scala 126:19]
  assign _GEN_110 = predicate_in_R_0_control == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_111 = _GEN_105 & _GEN_110; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_ready_R_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_ready_R_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_ready_R_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_ready_R_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  out_valid_R_8 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  out_valid_R_9 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  out_valid_R_10 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  out_valid_R_11 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  value = _RAND_24[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_25[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  state = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_4) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_5) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_6) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_6) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_6) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_7) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_7) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_7) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_8) begin
          out_ready_R_6 <= io_Out_6_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_6 <= 1'h0;
          end else begin
            if (_T_8) begin
              out_ready_R_6 <= io_Out_6_ready;
            end
          end
        end else begin
          if (_T_8) begin
            out_ready_R_6 <= io_Out_6_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_9) begin
          out_ready_R_7 <= io_Out_7_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_7 <= 1'h0;
          end else begin
            if (_T_9) begin
              out_ready_R_7 <= io_Out_7_ready;
            end
          end
        end else begin
          if (_T_9) begin
            out_ready_R_7 <= io_Out_7_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_8 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_10) begin
          out_ready_R_8 <= io_Out_8_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_8 <= 1'h0;
          end else begin
            if (_T_10) begin
              out_ready_R_8 <= io_Out_8_ready;
            end
          end
        end else begin
          if (_T_10) begin
            out_ready_R_8 <= io_Out_8_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_9 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_11) begin
          out_ready_R_9 <= io_Out_9_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_9 <= 1'h0;
          end else begin
            if (_T_11) begin
              out_ready_R_9 <= io_Out_9_ready;
            end
          end
        end else begin
          if (_T_11) begin
            out_ready_R_9 <= io_Out_9_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_10 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_12) begin
          out_ready_R_10 <= io_Out_10_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_10 <= 1'h0;
          end else begin
            if (_T_12) begin
              out_ready_R_10 <= io_Out_10_ready;
            end
          end
        end else begin
          if (_T_12) begin
            out_ready_R_10 <= io_Out_10_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_11 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_13) begin
          out_ready_R_11 <= io_Out_11_ready;
        end
      end else begin
        if (state) begin
          if (_T_38) begin
            out_ready_R_11 <= 1'h0;
          end else begin
            if (_T_13) begin
              out_ready_R_11 <= io_Out_11_ready;
            end
          end
        end else begin
          if (_T_13) begin
            out_ready_R_11 <= io_Out_11_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_0 <= _GEN_31;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_1 <= _GEN_32;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_2 <= _GEN_33;
      end else begin
        if (_T_4) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_3 <= _GEN_34;
      end else begin
        if (_T_5) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_4 <= _GEN_35;
      end else begin
        if (_T_6) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_5 <= _GEN_36;
      end else begin
        if (_T_7) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_6 <= _GEN_37;
      end else begin
        if (_T_8) begin
          out_valid_R_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_7 <= _GEN_38;
      end else begin
        if (_T_9) begin
          out_valid_R_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_8 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_8 <= _GEN_39;
      end else begin
        if (_T_10) begin
          out_valid_R_8 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_9 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_9 <= _GEN_40;
      end else begin
        if (_T_11) begin
          out_valid_R_9 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_10 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_10 <= _GEN_41;
      end else begin
        if (_T_12) begin
          out_valid_R_10 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_11 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_11 <= _GEN_42;
      end else begin
        if (_T_13) begin
          out_valid_R_11 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_17;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_21) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_21) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_21) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        predicate_valid_R_0 <= start;
      end else begin
        if (state) begin
          if (_T_38) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= start;
          end
        end else begin
          predicate_valid_R_0 <= start;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_24) begin
        state <= _GEN_44;
      end else begin
        if (state) begin
          if (_T_38) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_106 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup2615: Output fired @ %d, Mask: %d\n",predicate_in_R_0_taskID,value,predicate_control_R_0); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_111 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] bb_for_cond_cleanup2615: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_5(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_MaskBB_1_ready,
  output       io_MaskBB_1_valid,
  output [1:0] io_MaskBB_1_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output [4:0] io_Out_5_bits_taskID,
  output       io_Out_5_bits_control,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output [4:0] io_Out_6_bits_taskID,
  output       io_Out_6_bits_control,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output [4:0] io_Out_7_bits_taskID,
  output       io_Out_7_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_4;
  reg  out_ready_R_5; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_5;
  reg  out_ready_R_6; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_6;
  reg  out_ready_R_7; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_7;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_8;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_9;
  reg  out_valid_R_2; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_10;
  reg  out_valid_R_3; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_11;
  reg  out_valid_R_4; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_12;
  reg  out_valid_R_5; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_13;
  reg  out_valid_R_6; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_14;
  reg  out_valid_R_7; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_15;
  reg  mask_valid_R_0; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_16;
  reg  mask_valid_R_1; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_17;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 716:29]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[HandShaking.scala 716:29]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[HandShaking.scala 716:29]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[HandShaking.scala 716:29]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[HandShaking.scala 716:29]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[HandShaking.scala 716:29]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[HandShaking.scala 727:32]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[HandShaking.scala 727:32]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_18;
  wire [14:0] _T_14; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_19;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_20;
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_21;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_22;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_23;
  reg  predicate_control_R_1; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_24;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_25;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_26;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_27;
  wire  predicate; // @[BasicBlock.scala 75:58]
  wire [4:0] predicate_task; // @[BasicBlock.scala 76:62]
  wire  _T_19; // @[Decoupled.scala 40:37]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _T_21; // @[BasicBlock.scala 78:91]
  wire  _T_22; // @[BasicBlock.scala 78:91]
  wire  start; // @[BasicBlock.scala 78:107]
  wire [1:0] _T_27; // @[BasicBlock.scala 102:52]
  wire  _T_29; // @[Conditional.scala 37:30]
  wire  _GEN_29; // @[BasicBlock.scala 112:19]
  wire  _GEN_30; // @[BasicBlock.scala 112:19]
  wire  _GEN_31; // @[BasicBlock.scala 112:19]
  wire  _GEN_32; // @[BasicBlock.scala 112:19]
  wire  _GEN_33; // @[BasicBlock.scala 112:19]
  wire  _GEN_34; // @[BasicBlock.scala 112:19]
  wire  _GEN_35; // @[BasicBlock.scala 112:19]
  wire  _GEN_36; // @[BasicBlock.scala 112:19]
  wire  _GEN_37; // @[BasicBlock.scala 112:19]
  wire  _GEN_38; // @[BasicBlock.scala 112:19]
  wire  _GEN_39; // @[BasicBlock.scala 112:19]
  wire [7:0] _T_38; // @[HandShaking.scala 741:17]
  wire  _T_39; // @[HandShaking.scala 741:24]
  wire  _T_42; // @[BasicBlock.scala 126:19]
  wire  _T_43; // @[BasicBlock.scala 126:19]
  wire  _GEN_89; // @[BasicBlock.scala 126:19]
  wire  _GEN_90; // @[BasicBlock.scala 126:19]
  wire  _GEN_91; // @[BasicBlock.scala 126:19]
  wire  _GEN_92; // @[BasicBlock.scala 126:19]
  wire  _GEN_96; // @[BasicBlock.scala 132:19]
  wire  _GEN_97; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 716:29]
  assign _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 716:29]
  assign _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 716:29]
  assign _T_7 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_7 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 716:29]
  assign _T_8 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_8 ? 1'h0 : out_valid_R_6; // @[HandShaking.scala 716:29]
  assign _T_9 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_9 ? 1'h0 : out_valid_R_7; // @[HandShaking.scala 716:29]
  assign _T_10 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_10 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 727:32]
  assign _T_11 = io_MaskBB_1_ready & io_MaskBB_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_11 ? 1'h0 : mask_valid_R_1; // @[HandShaking.scala 727:32]
  assign _T_14 = value + 15'h1; // @[Counter.scala 38:22]
  assign predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 75:58]
  assign predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 76:62]
  assign _T_19 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _T_20 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _T_21 = _T_19 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_22 = _T_20 | predicate_valid_R_1; // @[BasicBlock.scala 78:91]
  assign start = _T_21 & _T_22; // @[BasicBlock.scala 78:107]
  assign _T_27 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:52]
  assign _T_29 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_29 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_30 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_31 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_32 = start | _GEN_7; // @[BasicBlock.scala 112:19]
  assign _GEN_33 = start | _GEN_9; // @[BasicBlock.scala 112:19]
  assign _GEN_34 = start | _GEN_11; // @[BasicBlock.scala 112:19]
  assign _GEN_35 = start | _GEN_13; // @[BasicBlock.scala 112:19]
  assign _GEN_36 = start | _GEN_15; // @[BasicBlock.scala 112:19]
  assign _GEN_37 = start | _GEN_17; // @[BasicBlock.scala 112:19]
  assign _GEN_38 = start | _GEN_19; // @[BasicBlock.scala 112:19]
  assign _GEN_39 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_38 = {out_ready_R_7,out_ready_R_6,out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_39 = _T_38 == 8'hff; // @[HandShaking.scala 741:24]
  assign _T_42 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_43 = _T_42 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 726:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_MaskBB_1_valid = mask_valid_R_1; // @[HandShaking.scala 726:24]
  assign io_MaskBB_1_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 715:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 715:21]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 715:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 715:21]
  assign io_Out_5_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_5_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 715:21]
  assign io_Out_6_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_6_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 715:21]
  assign io_Out_7_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_7_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 86:29]
  assign _GEN_89 = _T_29 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_90 = _GEN_89 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_91 = _GEN_90 & _T_39; // @[BasicBlock.scala 126:19]
  assign _GEN_92 = _GEN_91 & predicate; // @[BasicBlock.scala 126:19]
  assign _GEN_96 = predicate == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_97 = _GEN_91 & _GEN_96; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  mask_valid_R_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  value = _RAND_18[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  state = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_39) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_39) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_4) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_39) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_5) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_39) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_6) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_39) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_6) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_6) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_7) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_39) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_7) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_7) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_8) begin
          out_ready_R_6 <= io_Out_6_ready;
        end
      end else begin
        if (state) begin
          if (_T_39) begin
            out_ready_R_6 <= 1'h0;
          end else begin
            if (_T_8) begin
              out_ready_R_6 <= io_Out_6_ready;
            end
          end
        end else begin
          if (_T_8) begin
            out_ready_R_6 <= io_Out_6_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else begin
      if (_T_29) begin
        if (_T_9) begin
          out_ready_R_7 <= io_Out_7_ready;
        end
      end else begin
        if (state) begin
          if (_T_39) begin
            out_ready_R_7 <= 1'h0;
          end else begin
            if (_T_9) begin
              out_ready_R_7 <= io_Out_7_ready;
            end
          end
        end else begin
          if (_T_9) begin
            out_ready_R_7 <= io_Out_7_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_29) begin
        out_valid_R_0 <= _GEN_29;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_29) begin
        out_valid_R_1 <= _GEN_30;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_29) begin
        out_valid_R_2 <= _GEN_31;
      end else begin
        if (_T_4) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_29) begin
        out_valid_R_3 <= _GEN_32;
      end else begin
        if (_T_5) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_29) begin
        out_valid_R_4 <= _GEN_33;
      end else begin
        if (_T_6) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_29) begin
        out_valid_R_5 <= _GEN_34;
      end else begin
        if (_T_7) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else begin
      if (_T_29) begin
        out_valid_R_6 <= _GEN_35;
      end else begin
        if (_T_8) begin
          out_valid_R_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else begin
      if (_T_29) begin
        out_valid_R_7 <= _GEN_36;
      end else begin
        if (_T_9) begin
          out_valid_R_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_29) begin
        mask_valid_R_0 <= _GEN_37;
      end else begin
        if (_T_10) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_1 <= 1'h0;
    end else begin
      if (_T_29) begin
        mask_valid_R_1 <= _GEN_38;
      end else begin
        if (_T_11) begin
          mask_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_14;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_19) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_19) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_20) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_20) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_19) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_20) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_29) begin
        predicate_valid_R_0 <= _T_21;
      end else begin
        if (state) begin
          if (_T_39) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= _T_21;
          end
        end else begin
          predicate_valid_R_0 <= _T_21;
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_29) begin
        predicate_valid_R_1 <= _T_22;
      end else begin
        if (state) begin
          if (_T_39) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            predicate_valid_R_1 <= _T_22;
          end
        end else begin
          predicate_valid_R_1 <= _T_22;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_29) begin
        state <= _GEN_39;
      end else begin
        if (state) begin
          if (_T_39) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_92 & _T_43) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body2716: Output fired @ %d, Mask: %d\n",predicate_task,value,_T_27); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_97 & _T_43) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] bb_for_body2716: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_6(
  input        clock,
  input        reset,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output [4:0] io_Out_5_bits_taskID,
  output       io_Out_5_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_4;
  reg  out_ready_R_5; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_5;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_6;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_7;
  reg  out_valid_R_2; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_8;
  reg  out_valid_R_3; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_9;
  reg  out_valid_R_4; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_10;
  reg  out_valid_R_5; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_11;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 716:29]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[HandShaking.scala 716:29]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[HandShaking.scala 716:29]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[HandShaking.scala 716:29]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_12;
  wire [14:0] _T_11; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_13;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_14;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_15;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_16;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_17;
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  start; // @[BasicBlock.scala 78:91]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _GEN_19; // @[BasicBlock.scala 112:19]
  wire  _GEN_20; // @[BasicBlock.scala 112:19]
  wire  _GEN_21; // @[BasicBlock.scala 112:19]
  wire  _GEN_22; // @[BasicBlock.scala 112:19]
  wire  _GEN_23; // @[BasicBlock.scala 112:19]
  wire  _GEN_24; // @[BasicBlock.scala 112:19]
  wire  _GEN_26; // @[BasicBlock.scala 112:19]
  wire [5:0] _T_25; // @[HandShaking.scala 741:17]
  wire  _T_26; // @[HandShaking.scala 741:24]
  wire  _T_28; // @[BasicBlock.scala 126:19]
  wire  _T_29; // @[BasicBlock.scala 126:19]
  wire  _GEN_61; // @[BasicBlock.scala 126:19]
  wire  _GEN_62; // @[BasicBlock.scala 126:19]
  wire  _GEN_63; // @[BasicBlock.scala 126:19]
  wire  _GEN_64; // @[BasicBlock.scala 126:19]
  wire  _GEN_68; // @[BasicBlock.scala 132:19]
  wire  _GEN_69; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 716:29]
  assign _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 716:29]
  assign _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 716:29]
  assign _T_7 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_7 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 716:29]
  assign _T_11 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_15 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign start = _T_15 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_19 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_20 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_21 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_22 = start | _GEN_7; // @[BasicBlock.scala 112:19]
  assign _GEN_23 = start | _GEN_9; // @[BasicBlock.scala 112:19]
  assign _GEN_24 = start | _GEN_11; // @[BasicBlock.scala 112:19]
  assign _GEN_26 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_25 = {out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_26 = _T_25 == 6'h3f; // @[HandShaking.scala 741:24]
  assign _T_28 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_29 = _T_28 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 715:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 715:21]
  assign io_Out_3_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_3_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 715:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_4_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 715:21]
  assign io_Out_5_bits_taskID = predicate_in_R_0_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_5_bits_control = predicate_in_R_0_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign _GEN_61 = _T_18 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_62 = _GEN_61 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_63 = _GEN_62 & _T_26; // @[BasicBlock.scala 126:19]
  assign _GEN_64 = _GEN_63 & predicate_in_R_0_control; // @[BasicBlock.scala 126:19]
  assign _GEN_68 = predicate_in_R_0_control == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_69 = _GEN_63 & _GEN_68; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  value = _RAND_12[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_13[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  state = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_5) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_6) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_6) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_6) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_7) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_7) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_7) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        out_valid_R_0 <= _GEN_19;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        out_valid_R_1 <= _GEN_20;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_18) begin
        out_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_4) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_18) begin
        out_valid_R_3 <= _GEN_22;
      end else begin
        if (_T_5) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_18) begin
        out_valid_R_4 <= _GEN_23;
      end else begin
        if (_T_6) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_18) begin
        out_valid_R_5 <= _GEN_24;
      end else begin
        if (_T_7) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_11;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_15) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        predicate_valid_R_0 <= start;
      end else begin
        if (state) begin
          if (_T_26) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= start;
          end
        end else begin
          predicate_valid_R_0 <= start;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_26;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_64 & _T_29) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_cond_cleanup3317: Output fired @ %d, Mask: %d\n",predicate_in_R_0_taskID,value,predicate_control_R_0); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_69 & _T_29) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] bb_for_cond_cleanup3317: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_7(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_MaskBB_1_ready,
  output       io_MaskBB_1_valid,
  output [1:0] io_MaskBB_1_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output       io_Out_4_bits_control,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output [4:0] io_Out_5_bits_taskID,
  output       io_Out_5_bits_control,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output [4:0] io_Out_6_bits_taskID,
  output       io_Out_6_bits_control,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output [4:0] io_Out_7_bits_taskID,
  output       io_Out_7_bits_control,
  input        io_Out_8_ready,
  output       io_Out_8_valid,
  output [4:0] io_Out_8_bits_taskID,
  input        io_Out_9_ready,
  output       io_Out_9_valid,
  output [4:0] io_Out_9_bits_taskID,
  output       io_Out_9_bits_control,
  input        io_Out_10_ready,
  output       io_Out_10_valid,
  output [4:0] io_Out_10_bits_taskID,
  output       io_Out_10_bits_control,
  input        io_Out_11_ready,
  output       io_Out_11_valid,
  output [4:0] io_Out_11_bits_taskID,
  output       io_Out_11_bits_control,
  input        io_Out_12_ready,
  output       io_Out_12_valid,
  output [4:0] io_Out_12_bits_taskID,
  output       io_Out_12_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_4;
  reg  out_ready_R_5; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_5;
  reg  out_ready_R_6; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_6;
  reg  out_ready_R_7; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_7;
  reg  out_ready_R_8; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_8;
  reg  out_ready_R_9; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_9;
  reg  out_ready_R_10; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_10;
  reg  out_ready_R_11; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_11;
  reg  out_ready_R_12; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_12;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_13;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_14;
  reg  out_valid_R_2; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_15;
  reg  out_valid_R_3; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_16;
  reg  out_valid_R_4; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_17;
  reg  out_valid_R_5; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_18;
  reg  out_valid_R_6; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_19;
  reg  out_valid_R_7; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_20;
  reg  out_valid_R_8; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_21;
  reg  out_valid_R_9; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_22;
  reg  out_valid_R_10; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_23;
  reg  out_valid_R_11; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_24;
  reg  out_valid_R_12; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_25;
  reg  mask_valid_R_0; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_26;
  reg  mask_valid_R_1; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_27;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 716:29]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[HandShaking.scala 716:29]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[HandShaking.scala 716:29]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[HandShaking.scala 716:29]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[HandShaking.scala 716:29]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[HandShaking.scala 716:29]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[HandShaking.scala 716:29]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[HandShaking.scala 716:29]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[HandShaking.scala 716:29]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_23; // @[HandShaking.scala 716:29]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[HandShaking.scala 716:29]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_27; // @[HandShaking.scala 727:32]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[HandShaking.scala 727:32]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_28;
  wire [14:0] _T_19; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_29;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_30;
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_31;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_32;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_33;
  reg  predicate_control_R_1; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_34;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_35;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_36;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_37;
  wire  predicate; // @[BasicBlock.scala 75:58]
  wire [4:0] predicate_task; // @[BasicBlock.scala 76:62]
  wire  _T_24; // @[Decoupled.scala 40:37]
  wire  _T_25; // @[Decoupled.scala 40:37]
  wire  _T_26; // @[BasicBlock.scala 78:91]
  wire  _T_27; // @[BasicBlock.scala 78:91]
  wire  start; // @[BasicBlock.scala 78:107]
  wire [1:0] _T_32; // @[BasicBlock.scala 102:52]
  wire  _T_34; // @[Conditional.scala 37:30]
  wire  _GEN_39; // @[BasicBlock.scala 112:19]
  wire  _GEN_40; // @[BasicBlock.scala 112:19]
  wire  _GEN_41; // @[BasicBlock.scala 112:19]
  wire  _GEN_42; // @[BasicBlock.scala 112:19]
  wire  _GEN_43; // @[BasicBlock.scala 112:19]
  wire  _GEN_44; // @[BasicBlock.scala 112:19]
  wire  _GEN_45; // @[BasicBlock.scala 112:19]
  wire  _GEN_46; // @[BasicBlock.scala 112:19]
  wire  _GEN_47; // @[BasicBlock.scala 112:19]
  wire  _GEN_48; // @[BasicBlock.scala 112:19]
  wire  _GEN_49; // @[BasicBlock.scala 112:19]
  wire  _GEN_50; // @[BasicBlock.scala 112:19]
  wire  _GEN_51; // @[BasicBlock.scala 112:19]
  wire  _GEN_52; // @[BasicBlock.scala 112:19]
  wire  _GEN_53; // @[BasicBlock.scala 112:19]
  wire  _GEN_54; // @[BasicBlock.scala 112:19]
  wire [5:0] _T_41; // @[HandShaking.scala 741:17]
  wire [12:0] _T_48; // @[HandShaking.scala 741:17]
  wire  _T_49; // @[HandShaking.scala 741:24]
  wire  _T_52; // @[BasicBlock.scala 126:19]
  wire  _T_53; // @[BasicBlock.scala 126:19]
  wire  _GEN_124; // @[BasicBlock.scala 126:19]
  wire  _GEN_125; // @[BasicBlock.scala 126:19]
  wire  _GEN_126; // @[BasicBlock.scala 126:19]
  wire  _GEN_127; // @[BasicBlock.scala 126:19]
  wire  _GEN_131; // @[BasicBlock.scala 132:19]
  wire  _GEN_132; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 716:29]
  assign _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 716:29]
  assign _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 716:29]
  assign _T_7 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_7 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 716:29]
  assign _T_8 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_8 ? 1'h0 : out_valid_R_6; // @[HandShaking.scala 716:29]
  assign _T_9 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_9 ? 1'h0 : out_valid_R_7; // @[HandShaking.scala 716:29]
  assign _T_10 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_10 ? 1'h0 : out_valid_R_8; // @[HandShaking.scala 716:29]
  assign _T_11 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_11 ? 1'h0 : out_valid_R_9; // @[HandShaking.scala 716:29]
  assign _T_12 = io_Out_10_ready & io_Out_10_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_12 ? 1'h0 : out_valid_R_10; // @[HandShaking.scala 716:29]
  assign _T_13 = io_Out_11_ready & io_Out_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_23 = _T_13 ? 1'h0 : out_valid_R_11; // @[HandShaking.scala 716:29]
  assign _T_14 = io_Out_12_ready & io_Out_12_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_14 ? 1'h0 : out_valid_R_12; // @[HandShaking.scala 716:29]
  assign _T_15 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_27 = _T_15 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 727:32]
  assign _T_16 = io_MaskBB_1_ready & io_MaskBB_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_16 ? 1'h0 : mask_valid_R_1; // @[HandShaking.scala 727:32]
  assign _T_19 = value + 15'h1; // @[Counter.scala 38:22]
  assign predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 75:58]
  assign predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 76:62]
  assign _T_24 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _T_25 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _T_26 = _T_24 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_27 = _T_25 | predicate_valid_R_1; // @[BasicBlock.scala 78:91]
  assign start = _T_26 & _T_27; // @[BasicBlock.scala 78:107]
  assign _T_32 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:52]
  assign _T_34 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_39 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_40 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_41 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_42 = start | _GEN_7; // @[BasicBlock.scala 112:19]
  assign _GEN_43 = start | _GEN_9; // @[BasicBlock.scala 112:19]
  assign _GEN_44 = start | _GEN_11; // @[BasicBlock.scala 112:19]
  assign _GEN_45 = start | _GEN_13; // @[BasicBlock.scala 112:19]
  assign _GEN_46 = start | _GEN_15; // @[BasicBlock.scala 112:19]
  assign _GEN_47 = start | _GEN_17; // @[BasicBlock.scala 112:19]
  assign _GEN_48 = start | _GEN_19; // @[BasicBlock.scala 112:19]
  assign _GEN_49 = start | _GEN_21; // @[BasicBlock.scala 112:19]
  assign _GEN_50 = start | _GEN_23; // @[BasicBlock.scala 112:19]
  assign _GEN_51 = start | _GEN_25; // @[BasicBlock.scala 112:19]
  assign _GEN_52 = start | _GEN_27; // @[BasicBlock.scala 112:19]
  assign _GEN_53 = start | _GEN_29; // @[BasicBlock.scala 112:19]
  assign _GEN_54 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_41 = {out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_48 = {out_ready_R_12,out_ready_R_11,out_ready_R_10,out_ready_R_9,out_ready_R_8,out_ready_R_7,out_ready_R_6,_T_41}; // @[HandShaking.scala 741:17]
  assign _T_49 = _T_48 == 13'h1fff; // @[HandShaking.scala 741:24]
  assign _T_52 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_53 = _T_52 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 726:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_MaskBB_1_valid = mask_valid_R_1; // @[HandShaking.scala 726:24]
  assign io_MaskBB_1_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 715:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 715:21]
  assign io_Out_3_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 715:21]
  assign io_Out_4_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 715:21]
  assign io_Out_5_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_5_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 715:21]
  assign io_Out_6_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_6_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 715:21]
  assign io_Out_7_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_7_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_8_valid = out_valid_R_8; // @[HandShaking.scala 715:21]
  assign io_Out_8_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_9_valid = out_valid_R_9; // @[HandShaking.scala 715:21]
  assign io_Out_9_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_9_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_10_valid = out_valid_R_10; // @[HandShaking.scala 715:21]
  assign io_Out_10_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_10_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_11_valid = out_valid_R_11; // @[HandShaking.scala 715:21]
  assign io_Out_11_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_11_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_12_valid = out_valid_R_12; // @[HandShaking.scala 715:21]
  assign io_Out_12_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_12_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 86:29]
  assign _GEN_124 = _T_34 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_125 = _GEN_124 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_126 = _GEN_125 & _T_49; // @[BasicBlock.scala 126:19]
  assign _GEN_127 = _GEN_126 & predicate; // @[BasicBlock.scala 126:19]
  assign _GEN_131 = predicate == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_132 = _GEN_126 & _GEN_131; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_ready_R_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_ready_R_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_ready_R_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_ready_R_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_ready_R_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  out_valid_R_8 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  out_valid_R_9 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  out_valid_R_10 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  out_valid_R_11 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  out_valid_R_12 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mask_valid_R_1 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  value = _RAND_28[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_29[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  state = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_4) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_5) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_6) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_6) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_6) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_7) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_7) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_7) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_8) begin
          out_ready_R_6 <= io_Out_6_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_6 <= 1'h0;
          end else begin
            if (_T_8) begin
              out_ready_R_6 <= io_Out_6_ready;
            end
          end
        end else begin
          if (_T_8) begin
            out_ready_R_6 <= io_Out_6_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_9) begin
          out_ready_R_7 <= io_Out_7_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_7 <= 1'h0;
          end else begin
            if (_T_9) begin
              out_ready_R_7 <= io_Out_7_ready;
            end
          end
        end else begin
          if (_T_9) begin
            out_ready_R_7 <= io_Out_7_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_8 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_10) begin
          out_ready_R_8 <= io_Out_8_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_8 <= 1'h0;
          end else begin
            if (_T_10) begin
              out_ready_R_8 <= io_Out_8_ready;
            end
          end
        end else begin
          if (_T_10) begin
            out_ready_R_8 <= io_Out_8_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_9 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_11) begin
          out_ready_R_9 <= io_Out_9_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_9 <= 1'h0;
          end else begin
            if (_T_11) begin
              out_ready_R_9 <= io_Out_9_ready;
            end
          end
        end else begin
          if (_T_11) begin
            out_ready_R_9 <= io_Out_9_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_10 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_12) begin
          out_ready_R_10 <= io_Out_10_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_10 <= 1'h0;
          end else begin
            if (_T_12) begin
              out_ready_R_10 <= io_Out_10_ready;
            end
          end
        end else begin
          if (_T_12) begin
            out_ready_R_10 <= io_Out_10_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_11 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_13) begin
          out_ready_R_11 <= io_Out_11_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_11 <= 1'h0;
          end else begin
            if (_T_13) begin
              out_ready_R_11 <= io_Out_11_ready;
            end
          end
        end else begin
          if (_T_13) begin
            out_ready_R_11 <= io_Out_11_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_12 <= 1'h0;
    end else begin
      if (_T_34) begin
        if (_T_14) begin
          out_ready_R_12 <= io_Out_12_ready;
        end
      end else begin
        if (state) begin
          if (_T_49) begin
            out_ready_R_12 <= 1'h0;
          end else begin
            if (_T_14) begin
              out_ready_R_12 <= io_Out_12_ready;
            end
          end
        end else begin
          if (_T_14) begin
            out_ready_R_12 <= io_Out_12_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_0 <= _GEN_39;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_1 <= _GEN_40;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_2 <= _GEN_41;
      end else begin
        if (_T_4) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_3 <= _GEN_42;
      end else begin
        if (_T_5) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_4 <= _GEN_43;
      end else begin
        if (_T_6) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_5 <= _GEN_44;
      end else begin
        if (_T_7) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_6 <= _GEN_45;
      end else begin
        if (_T_8) begin
          out_valid_R_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_7 <= _GEN_46;
      end else begin
        if (_T_9) begin
          out_valid_R_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_8 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_8 <= _GEN_47;
      end else begin
        if (_T_10) begin
          out_valid_R_8 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_9 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_9 <= _GEN_48;
      end else begin
        if (_T_11) begin
          out_valid_R_9 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_10 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_10 <= _GEN_49;
      end else begin
        if (_T_12) begin
          out_valid_R_10 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_11 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_11 <= _GEN_50;
      end else begin
        if (_T_13) begin
          out_valid_R_11 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_12 <= 1'h0;
    end else begin
      if (_T_34) begin
        out_valid_R_12 <= _GEN_51;
      end else begin
        if (_T_14) begin
          out_valid_R_12 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_34) begin
        mask_valid_R_0 <= _GEN_52;
      end else begin
        if (_T_15) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_1 <= 1'h0;
    end else begin
      if (_T_34) begin
        mask_valid_R_1 <= _GEN_53;
      end else begin
        if (_T_16) begin
          mask_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_19;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_24) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_24) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_25) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_25) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_25) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_34) begin
        predicate_valid_R_0 <= _T_26;
      end else begin
        if (state) begin
          if (_T_49) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= _T_26;
          end
        end else begin
          predicate_valid_R_0 <= _T_26;
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_34) begin
        predicate_valid_R_1 <= _T_27;
      end else begin
        if (state) begin
          if (_T_49) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            predicate_valid_R_1 <= _T_27;
          end
        end else begin
          predicate_valid_R_1 <= _T_27;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_34) begin
        state <= _GEN_54;
      end else begin
        if (state) begin
          if (_T_49) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & _T_53) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [BB]   bb_for_body3418: Output fired @ %d, Mask: %d\n",predicate_task,value,_T_32); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_132 & _T_53) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] bb_for_body3418: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  assign io_out = io_in1 + io_in2; // @[Alu.scala 237:10]
endmodule
module ComputeNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add0: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_1(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire  _T_20; // @[Alu.scala 190:38]
  assign _T_20 = io_in1 > io_in2; // @[Alu.scala 190:38]
  assign io_out = {{31'd0}, _T_20}; // @[Alu.scala 237:10]
endmodule
module ComputeNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] icmp_cmp1421: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output [4:0]  io_TrueOutput_0_bits_taskID,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg [4:0] output_true_R_taskID; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_8;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_9;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_10;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_12;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_13;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_14;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_15;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_taskID = output_true_R_taskID; // @[BranchNode.scala 1259:27]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_R_control = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_R_control = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_true_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_taskID <= 5'h0;
          end else begin
            output_true_R_taskID <= task_id;
          end
        end else begin
          output_true_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_2: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_2: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add43: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] icmp_cmp51394: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add125: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] icmp_cmp131376: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_7: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_7: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_1(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_8: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_8: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module RetNode2(
  input        clock,
  input        reset,
  output       io_In_enable_ready,
  input        io_In_enable_valid,
  input  [4:0] io_In_enable_bits_taskID,
  input        io_In_enable_bits_control,
  input        io_Out_ready,
  output       io_Out_valid,
  output [4:0] io_Out_bits_enable_taskID,
  output       io_Out_bits_enable_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg  state; // @[RetNode.scala 131:22]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[RetNode.scala 134:31]
  reg [31:0] _RAND_2;
  reg [4:0] output_R_enable_taskID; // @[RetNode.scala 140:25]
  reg [31:0] _RAND_3;
  reg  output_R_enable_control; // @[RetNode.scala 140:25]
  reg [31:0] _RAND_4;
  reg  out_ready_R; // @[RetNode.scala 141:28]
  reg [31:0] _RAND_5;
  reg  out_valid_R; // @[RetNode.scala 142:28]
  reg [31:0] _RAND_6;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[RetNode.scala 172:23]
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _GEN_8; // @[RetNode.scala 179:28]
  wire  _GEN_9; // @[RetNode.scala 179:28]
  wire  _T_13; // @[RetNode.scala 198:17]
  wire  _T_14; // @[RetNode.scala 198:17]
  wire  _GEN_22; // @[RetNode.scala 198:17]
  wire  _GEN_23; // @[RetNode.scala 198:17]
  wire  _GEN_24; // @[RetNode.scala 198:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_9 = io_In_enable_ready & io_In_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_10 ? 1'h0 : out_valid_R; // @[RetNode.scala 172:23]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_8 = enable_valid_R | _GEN_5; // @[RetNode.scala 179:28]
  assign _GEN_9 = enable_valid_R | state; // @[RetNode.scala 179:28]
  assign _T_13 = $unsigned(reset); // @[RetNode.scala 198:17]
  assign _T_14 = _T_13 == 1'h0; // @[RetNode.scala 198:17]
  assign io_In_enable_ready = ~ enable_valid_R; // @[RetNode.scala 153:22]
  assign io_Out_valid = out_valid_R; // @[RetNode.scala 170:16]
  assign io_Out_bits_enable_taskID = output_R_enable_taskID; // @[RetNode.scala 169:15]
  assign io_Out_bits_enable_control = output_R_enable_control; // @[RetNode.scala 169:15]
  assign _GEN_22 = _T_11 == 1'h0; // @[RetNode.scala 198:17]
  assign _GEN_23 = _GEN_22 & state; // @[RetNode.scala 198:17]
  assign _GEN_24 = _GEN_23 & out_ready_R; // @[RetNode.scala 198:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  output_R_enable_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_enable_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_9;
      end else begin
        if (state) begin
          if (out_ready_R) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_9) begin
          enable_valid_R <= io_In_enable_valid;
        end
      end else begin
        if (state) begin
          if (out_ready_R) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_9) begin
              enable_valid_R <= io_In_enable_valid;
            end
          end
        end else begin
          if (_T_9) begin
            enable_valid_R <= io_In_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      output_R_enable_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        output_R_enable_taskID <= io_In_enable_bits_taskID;
      end
    end
    if (reset) begin
      output_R_enable_control <= 1'h0;
    end else begin
      if (_T_9) begin
        output_R_enable_control <= io_In_enable_bits_control;
      end
    end
    if (reset) begin
      out_ready_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_10) begin
          out_ready_R <= io_Out_ready;
        end
      end else begin
        if (state) begin
          if (out_ready_R) begin
            out_ready_R <= 1'h0;
          end else begin
            if (_T_10) begin
              out_ready_R <= io_Out_ready;
            end
          end
        end else begin
          if (_T_10) begin
            out_ready_R <= io_Out_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        out_valid_R <= _GEN_8;
      end else begin
        if (state) begin
          if (out_ready_R) begin
            out_valid_R <= 1'h0;
          end else begin
            if (_T_10) begin
              out_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            out_valid_R <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_24 & _T_14) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [RET] ret_9: Output fired @ %d\n",output_R_enable_taskID,value); // @[RetNode.scala 198:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  input  [31:0] io_InData_0_bits_data,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_0_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_6;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_7;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_8;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_9;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_10;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_11;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_12;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_17; // @[Bitwise.scala 108:18]
  wire  _T_18; // @[Bitwise.scala 108:44]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_13;
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _T_25; // @[PhiNode.scala 268:37]
  wire  _T_26; // @[PhiNode.scala 277:27]
  wire  _T_27; // @[PhiNode.scala 283:19]
  wire  _T_28; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_32; // @[PhiNode.scala 283:19]
  wire  _GEN_35; // @[PhiNode.scala 277:46]
  wire  _GEN_36; // @[PhiNode.scala 277:46]
  wire  _T_31; // @[Conditional.scala 37:30]
  wire  _T_32; // @[PhiNode.scala 299:31]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_70; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_108; // @[Conditional.scala 39:67]
  wire  _GEN_138; // @[PhiNode.scala 283:19]
  wire  _GEN_139; // @[PhiNode.scala 283:19]
  wire  _GEN_141; // @[PhiNode.scala 291:19]
  wire  _GEN_142; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_17 = mask_R[0]; // @[Bitwise.scala 108:18]
  assign _T_18 = mask_R[1]; // @[Bitwise.scala 108:44]
  assign _T_19 = {_T_17,_T_18}; // @[Cat.scala 29:58]
  assign sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  assign _GEN_19 = sel ? in_data_R_1_data : in_data_R_0_data; // @[PhiNode.scala 253:20]
  assign _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_20 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = _T_21 | fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 265:74]
  assign _T_24 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_25 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_26 = enable_valid_R & _T_25; // @[PhiNode.scala 277:27]
  assign _T_27 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_28 = _T_27 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_32 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_35 = _T_26 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_36 = _T_26 | _GEN_23; // @[PhiNode.scala 277:46]
  assign _T_31 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_32 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_70 = _T_36 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_108 = _T_31 ? _GEN_19 : _GEN_70; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_24 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_data = _T_24 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_138 = _T_24 & _T_26; // @[PhiNode.scala 283:19]
  assign _GEN_139 = _GEN_138 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_141 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_142 = _GEN_138 & _GEN_141; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mask_R = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mask_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  fire_R_0 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fire_R_1 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  state = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_data <= 32'h0;
    end else begin
      if (_T_24) begin
        if (_T_14) begin
          in_data_R_0_data <= io_InData_0_bits_data;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_R_0_data <= 32'h0;
          end else begin
            if (_T_14) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_R_0_data <= 32'h0;
            end else begin
              if (_T_14) begin
                in_data_R_0_data <= io_InData_0_bits_data;
              end
            end
          end else begin
            if (_T_14) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_24) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_24) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_0 <= _GEN_35;
      end else begin
        if (_T_20) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_1 <= _GEN_36;
      end else begin
        if (_T_21) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        fire_R_1 <= _GEN_22;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            fire_R_1 <= 1'h0;
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_1 <= 1'h0;
            end else begin
              fire_R_1 <= _GEN_22;
            end
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_139 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_pw_conv_reduction_s1_k_014310: Output fired @ %d, Value: %d\n",_GEN_32,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_142 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_pw_conv_reduction_s1_k_014310: Output flushed @ %d, Value: %d\n",_GEN_32,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_6(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  assign io_out = io_in1 - io_in2; // @[Alu.scala 237:10]
endmodule
module ComputeNode_6(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_6 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_sub11: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_7(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire [63:0] _T_24; // @[Alu.scala 196:32]
  assign _T_24 = io_in1 * io_in2; // @[Alu.scala 196:32]
  assign io_out = _T_24[31:0]; // @[Alu.scala 237:10]
endmodule
module ComputeNode_7(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_7 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_mul112: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output [4:0]  io_TrueOutput_0_bits_taskID,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg [4:0] output_true_R_taskID; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_8;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_9;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_10;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_12;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_13;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_14;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_15;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_taskID = output_true_R_taskID; // @[BranchNode.scala 1259:27]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_R_control = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_R_control = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_true_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_taskID <= 5'h0;
          end else begin
            output_true_R_taskID <= task_id;
          end
        end else begin
          output_true_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_13: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_13: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_2(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_14: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_14: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_3(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_15: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_15: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_8(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_inc6416: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_9(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire  _T_21; // @[Alu.scala 191:38]
  assign _T_21 = io_in1 == io_in2; // @[Alu.scala 191:38]
  assign io_out = {{31'd0}, _T_21}; // @[Alu.scala 237:10]
endmodule
module ComputeNode_9(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_9 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] icmp_exitcond14817: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_8;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_9;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_10;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_12;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_13;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_14;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_18: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_18: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  input  [31:0] io_InData_0_bits_data,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [31:0] io_Out_2_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_0_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_6;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_7;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_8;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_9;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_10;
  reg  out_valid_R_2; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_11;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_12;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_13;
  reg  fire_R_2; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_14;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_17; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  _T_19; // @[Decoupled.scala 40:37]
  wire  _GEN_24; // @[PhiNode.scala 258:26]
  wire  _GEN_25; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  wire  fire_mask_2; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_15;
  wire  _T_23; // @[Conditional.scala 37:30]
  wire  _T_24; // @[PhiNode.scala 268:37]
  wire  _T_25; // @[PhiNode.scala 277:27]
  wire  _T_26; // @[PhiNode.scala 283:19]
  wire  _T_27; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_34; // @[PhiNode.scala 283:19]
  wire  _GEN_37; // @[PhiNode.scala 277:46]
  wire  _GEN_38; // @[PhiNode.scala 277:46]
  wire  _GEN_39; // @[PhiNode.scala 277:46]
  wire  _T_30; // @[Conditional.scala 37:30]
  wire  _T_31; // @[PhiNode.scala 299:31]
  wire  _T_32; // @[PhiNode.scala 299:31]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_75; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_118; // @[Conditional.scala 39:67]
  wire  _GEN_156; // @[PhiNode.scala 283:19]
  wire  _GEN_157; // @[PhiNode.scala 283:19]
  wire  _GEN_159; // @[PhiNode.scala 291:19]
  wire  _GEN_160; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign sel = mask_R[1]; // @[CircuitMath.scala 30:8]
  assign _GEN_19 = sel ? in_data_R_1_data : in_data_R_0_data; // @[PhiNode.scala 253:20]
  assign _T_17 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_17 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_17 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_18 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = _T_18 | fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_18 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign _T_19 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_24 = _T_19 | fire_R_2; // @[PhiNode.scala 258:26]
  assign _GEN_25 = _T_19 ? 1'h0 : out_valid_R_2; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_17; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_18; // @[PhiNode.scala 265:74]
  assign fire_mask_2 = fire_R_2 | _T_19; // @[PhiNode.scala 265:74]
  assign _T_23 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_24 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_25 = enable_valid_R & _T_24; // @[PhiNode.scala 277:27]
  assign _T_26 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_27 = _T_26 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_34 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_37 = _T_25 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_38 = _T_25 | _GEN_23; // @[PhiNode.scala 277:46]
  assign _GEN_39 = _T_25 | _GEN_25; // @[PhiNode.scala 277:46]
  assign _T_30 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_31 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_32 = _T_31 & fire_mask_2; // @[PhiNode.scala 299:31]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_75 = _T_36 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_118 = _T_30 ? _GEN_19 : _GEN_75; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_23 ? _GEN_19 : _GEN_118; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_data = _T_23 ? _GEN_19 : _GEN_118; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_2_valid = out_valid_R_2; // @[PhiNode.scala 254:21]
  assign io_Out_2_bits_data = _T_23 ? _GEN_19 : _GEN_118; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_156 = _T_23 & _T_25; // @[PhiNode.scala 283:19]
  assign _GEN_157 = _GEN_156 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_159 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_160 = _GEN_156 & _GEN_159; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mask_R = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mask_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fire_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_R_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_R_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_data <= 32'h0;
    end else begin
      if (_T_23) begin
        if (_T_14) begin
          in_data_R_0_data <= io_InData_0_bits_data;
        end
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            in_data_R_0_data <= 32'h0;
          end else begin
            if (_T_14) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_R_0_data <= 32'h0;
            end else begin
              if (_T_14) begin
                in_data_R_0_data <= io_InData_0_bits_data;
              end
            end
          end else begin
            if (_T_14) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_23) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_23) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_23) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_23) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_23) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_23) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_23) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_23) begin
        out_valid_R_0 <= _GEN_37;
      end else begin
        if (_T_17) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_23) begin
        out_valid_R_1 <= _GEN_38;
      end else begin
        if (_T_18) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_23) begin
        out_valid_R_2 <= _GEN_39;
      end else begin
        if (_T_19) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_23) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_23) begin
        fire_R_1 <= _GEN_22;
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            fire_R_1 <= 1'h0;
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_1 <= 1'h0;
            end else begin
              fire_R_1 <= _GEN_22;
            end
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end
      end
    end
    if (reset) begin
      fire_R_2 <= 1'h0;
    end else begin
      if (_T_23) begin
        fire_R_2 <= _GEN_24;
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            fire_R_2 <= 1'h0;
          end else begin
            fire_R_2 <= _GEN_24;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_2 <= 1'h0;
            end else begin
              fire_R_2 <= _GEN_24;
            end
          end else begin
            fire_R_2 <= _GEN_24;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_23) begin
        if (_T_25) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_30) begin
          if (_T_32) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_27) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_pw_conv_reduction_s1_y_014019: Output fired @ %d, Value: %d\n",_GEN_34,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_27) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_pw_conv_reduction_s1_y_014019: Output flushed @ %d, Value: %d\n",_GEN_34,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output [4:0]  io_TrueOutput_0_bits_taskID,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg [4:0] output_true_R_taskID; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_8;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_9;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_10;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_12;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_13;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_14;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_15;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_taskID = output_true_R_taskID; // @[BranchNode.scala 1259:27]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_R_control = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_R_control = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_true_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_taskID <= 5'h0;
          end else begin
            output_true_R_taskID <= task_id;
          end
        end else begin
          output_true_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_20: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_20: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_10(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_6 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_sub821: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_11(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_reass_add22: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_12(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_7 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_reass_mul23: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_4(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_24: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_24: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_5(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_25: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_25: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_13(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_inc6126: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_14(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_9 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] icmp_exitcond14727: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_8;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_9;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_10;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_12;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_13;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_14;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_28: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_28: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  input  [31:0] io_InData_0_bits_data,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [31:0] io_Out_2_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_0_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_6;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_7;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_8;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_9;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_10;
  reg  out_valid_R_2; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_11;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_12;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_13;
  reg  fire_R_2; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_14;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_17; // @[Bitwise.scala 108:18]
  wire  _T_18; // @[Bitwise.scala 108:44]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  _T_22; // @[Decoupled.scala 40:37]
  wire  _GEN_24; // @[PhiNode.scala 258:26]
  wire  _GEN_25; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  wire  fire_mask_2; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_15;
  wire  _T_26; // @[Conditional.scala 37:30]
  wire  _T_27; // @[PhiNode.scala 268:37]
  wire  _T_28; // @[PhiNode.scala 277:27]
  wire  _T_29; // @[PhiNode.scala 283:19]
  wire  _T_30; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_34; // @[PhiNode.scala 283:19]
  wire  _GEN_37; // @[PhiNode.scala 277:46]
  wire  _GEN_38; // @[PhiNode.scala 277:46]
  wire  _GEN_39; // @[PhiNode.scala 277:46]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_34; // @[PhiNode.scala 299:31]
  wire  _T_35; // @[PhiNode.scala 299:31]
  wire  _T_39; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_75; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_118; // @[Conditional.scala 39:67]
  wire  _GEN_156; // @[PhiNode.scala 283:19]
  wire  _GEN_157; // @[PhiNode.scala 283:19]
  wire  _GEN_159; // @[PhiNode.scala 291:19]
  wire  _GEN_160; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_17 = mask_R[0]; // @[Bitwise.scala 108:18]
  assign _T_18 = mask_R[1]; // @[Bitwise.scala 108:44]
  assign _T_19 = {_T_17,_T_18}; // @[Cat.scala 29:58]
  assign sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  assign _GEN_19 = sel ? in_data_R_1_data : in_data_R_0_data; // @[PhiNode.scala 253:20]
  assign _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_20 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = _T_21 | fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign _T_22 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_24 = _T_22 | fire_R_2; // @[PhiNode.scala 258:26]
  assign _GEN_25 = _T_22 ? 1'h0 : out_valid_R_2; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 265:74]
  assign fire_mask_2 = fire_R_2 | _T_22; // @[PhiNode.scala 265:74]
  assign _T_26 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_27 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_28 = enable_valid_R & _T_27; // @[PhiNode.scala 277:27]
  assign _T_29 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_30 = _T_29 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_34 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_37 = _T_28 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_38 = _T_28 | _GEN_23; // @[PhiNode.scala 277:46]
  assign _GEN_39 = _T_28 | _GEN_25; // @[PhiNode.scala 277:46]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_34 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_35 = _T_34 & fire_mask_2; // @[PhiNode.scala 299:31]
  assign _T_39 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_75 = _T_39 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_118 = _T_33 ? _GEN_19 : _GEN_75; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_26 ? _GEN_19 : _GEN_118; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_data = _T_26 ? _GEN_19 : _GEN_118; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_2_valid = out_valid_R_2; // @[PhiNode.scala 254:21]
  assign io_Out_2_bits_data = _T_26 ? _GEN_19 : _GEN_118; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_156 = _T_26 & _T_28; // @[PhiNode.scala 283:19]
  assign _GEN_157 = _GEN_156 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_159 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_160 = _GEN_156 & _GEN_159; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mask_R = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mask_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fire_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_R_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_R_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_data <= 32'h0;
    end else begin
      if (_T_26) begin
        if (_T_14) begin
          in_data_R_0_data <= io_InData_0_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            in_data_R_0_data <= 32'h0;
          end else begin
            if (_T_14) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              in_data_R_0_data <= 32'h0;
            end else begin
              if (_T_14) begin
                in_data_R_0_data <= io_InData_0_bits_data;
              end
            end
          end else begin
            if (_T_14) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_26) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_26) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_26) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_26) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_26) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_26) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_26) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_26) begin
        out_valid_R_0 <= _GEN_37;
      end else begin
        if (_T_20) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_26) begin
        out_valid_R_1 <= _GEN_38;
      end else begin
        if (_T_21) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_26) begin
        out_valid_R_2 <= _GEN_39;
      end else begin
        if (_T_22) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_26) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_26) begin
        fire_R_1 <= _GEN_22;
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            fire_R_1 <= 1'h0;
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              fire_R_1 <= 1'h0;
            end else begin
              fire_R_1 <= _GEN_22;
            end
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end
      end
    end
    if (reset) begin
      fire_R_2 <= 1'h0;
    end else begin
      if (_T_26) begin
        fire_R_2 <= _GEN_24;
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            fire_R_2 <= 1'h0;
          end else begin
            fire_R_2 <= _GEN_24;
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              fire_R_2 <= 1'h0;
            end else begin
              fire_R_2 <= _GEN_24;
            end
          end else begin
            fire_R_2 <= _GEN_24;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_26) begin
        if (_T_28) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_33) begin
          if (_T_35) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_39) begin
            if (_T_35) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_157 & _T_30) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_pw_conv_reduction_s1_x_013829: Output fired @ %d, Value: %d\n",_GEN_34,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_160 & _T_30) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_pw_conv_reduction_s1_x_013829: Output flushed @ %d, Value: %d\n",_GEN_34,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_15(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_6 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_sub1630: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_16(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_6 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add1031: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_17(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add1732: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [GEP] Gep_arrayidx5033: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_6(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_34: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_34: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_18(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_inc5835: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_19(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_9 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] icmp_exitcond14636: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_8;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_9;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_10;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_12;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_13;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_14;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_37: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_37: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_4;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_5;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_6;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_7;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_8;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_9;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_10;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_11;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_17; // @[Bitwise.scala 108:18]
  wire  _T_18; // @[Bitwise.scala 108:44]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_12;
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _T_25; // @[PhiNode.scala 268:37]
  wire  _T_26; // @[PhiNode.scala 277:27]
  wire  _T_27; // @[PhiNode.scala 283:19]
  wire  _T_28; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_32; // @[PhiNode.scala 283:19]
  wire  _GEN_35; // @[PhiNode.scala 277:46]
  wire  _GEN_36; // @[PhiNode.scala 277:46]
  wire  _T_31; // @[Conditional.scala 37:30]
  wire  _T_32; // @[PhiNode.scala 299:31]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_70; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_108; // @[Conditional.scala 39:67]
  wire  _GEN_138; // @[PhiNode.scala 283:19]
  wire  _GEN_139; // @[PhiNode.scala 283:19]
  wire  _GEN_141; // @[PhiNode.scala 291:19]
  wire  _GEN_142; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_17 = mask_R[0]; // @[Bitwise.scala 108:18]
  assign _T_18 = mask_R[1]; // @[Bitwise.scala 108:44]
  assign _T_19 = {_T_17,_T_18}; // @[Cat.scala 29:58]
  assign sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  assign _GEN_19 = sel ? in_data_R_1_data : 32'h0; // @[PhiNode.scala 253:20]
  assign _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_20 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = _T_21 | fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 265:74]
  assign _T_24 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_25 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_26 = enable_valid_R & _T_25; // @[PhiNode.scala 277:27]
  assign _T_27 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_28 = _T_27 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_32 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_35 = _T_26 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_36 = _T_26 | _GEN_23; // @[PhiNode.scala 277:46]
  assign _T_31 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_32 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_70 = _T_36 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_108 = _T_31 ? _GEN_19 : _GEN_70; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_24 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_data = _T_24 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_138 = _T_24 & _T_26; // @[PhiNode.scala 283:19]
  assign _GEN_139 = _GEN_138 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_141 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_142 = _GEN_138 & _GEN_141; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mask_R = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mask_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fire_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  fire_R_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_24) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_24) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_0 <= _GEN_35;
      end else begin
        if (_T_20) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_1 <= _GEN_36;
      end else begin
        if (_T_21) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        fire_R_1 <= _GEN_22;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            fire_R_1 <= 1'h0;
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_1 <= 1'h0;
            end else begin
              fire_R_1 <= _GEN_22;
            end
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_139 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_pw_conv_reduction_s1_r_pw__x_013638: Output fired @ %d, Value: %d\n",_GEN_32,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_142 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_pw_conv_reduction_s1_r_pw__x_013638: Output flushed @ %d, Value: %d\n",_GEN_32,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_20(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_7 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_mul2239: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_21(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add2340: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_7(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_41: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_41: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  input  [31:0] io_InData_0_bits_data,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_0_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_2;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_10; // @[PhiNode.scala 258:26]
  wire  _GEN_11; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_7;
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[PhiNode.scala 277:27]
  wire  _T_18; // @[PhiNode.scala 283:19]
  wire  _T_19; // @[PhiNode.scala 283:19]
  wire  _GEN_13; // @[PhiNode.scala 277:46]
  wire  _T_22; // @[Conditional.scala 37:30]
  wire  _T_25; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_31; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_56; // @[Conditional.scala 39:67]
  wire  _GEN_74; // @[PhiNode.scala 283:19]
  wire  _GEN_75; // @[PhiNode.scala 283:19]
  wire  _GEN_77; // @[PhiNode.scala 291:19]
  wire  _GEN_78; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_11 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_13 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_13 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_14 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_10 = _T_14 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_11 = _T_14 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_14; // @[PhiNode.scala 265:74]
  assign _T_16 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & in_data_valid_R_0; // @[PhiNode.scala 277:27]
  assign _T_18 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_19 = _T_18 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_13 = _T_17 | _GEN_11; // @[PhiNode.scala 277:46]
  assign _T_22 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_25 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_31 = _T_25 ? 32'h0 : in_data_R_0_data; // @[Conditional.scala 39:67]
  assign _GEN_56 = _T_22 ? in_data_R_0_data : _GEN_31; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_16 ? in_data_R_0_data : _GEN_56; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_74 = _T_16 & _T_17; // @[PhiNode.scala 283:19]
  assign _GEN_75 = _GEN_74 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_77 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_78 = _GEN_74 & _GEN_77; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_control = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_data <= 32'h0;
    end else begin
      if (_T_16) begin
        if (_T_13) begin
          in_data_R_0_data <= io_InData_0_bits_data;
        end
      end else begin
        if (_T_22) begin
          if (fire_mask_0) begin
            in_data_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end else begin
          if (_T_25) begin
            if (fire_mask_0) begin
              in_data_R_0_data <= 32'h0;
            end else begin
              if (_T_13) begin
                in_data_R_0_data <= io_InData_0_bits_data;
              end
            end
          end else begin
            if (_T_13) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_22) begin
          if (fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_25) begin
            if (fire_mask_0) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_11) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_22) begin
          if (fire_mask_0) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_11) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_25) begin
            if (fire_mask_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_11) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_11) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_22) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_25) begin
            if (fire_mask_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        out_valid_R_0 <= _GEN_13;
      end else begin
        if (_T_14) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        fire_R_0 <= _GEN_10;
      end else begin
        if (_T_22) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_10;
          end
        end else begin
          if (_T_25) begin
            if (fire_mask_0) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_10;
            end
          end else begin
            fire_R_0 <= _GEN_10;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_16) begin
        if (_T_17) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_22) begin
          if (fire_mask_0) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_25) begin
            if (fire_mask_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phiadd38_lcssa_lcssa42: Output fired @ %d, Value: %d\n",io_InData_0_bits_taskID,value,in_data_R_0_data); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_78 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phiadd38_lcssa_lcssa42: Output flushed @ %d, Value: %d\n",io_InData_0_bits_taskID,value,in_data_R_0_data); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_22(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_7 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h3;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_mul4443: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SextNode(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[SextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[SextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[SextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[SextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[SextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[SextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[SextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[SextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[SextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[SextNode.scala 84:26]
  wire  _GEN_9; // @[SextNode.scala 84:26]
  wire  fire_mask_0; // @[SextNode.scala 90:74]
  reg  state; // @[SextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[SextNode.scala 93:27]
  wire  _T_16; // @[SextNode.scala 97:26]
  wire  _T_17; // @[SextNode.scala 110:28]
  wire  _T_18; // @[SextNode.scala 117:17]
  wire  _T_19; // @[SextNode.scala 117:17]
  wire  _GEN_10; // @[SextNode.scala 110:47]
  wire  _GEN_11; // @[SextNode.scala 110:47]
  wire  _GEN_42; // @[SextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[SextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[SextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[SextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[SextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[SextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[SextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[SextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[SextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[SextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[SextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[SextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[SextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[SextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[SextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[SextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[SextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[SextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[SextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] sextconv4744: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[SextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOAD] ld_45: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOAD] ld_45: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOAD] ld_45: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_23(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add5246: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [STORE]st_47: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_24(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_inc5548: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_25(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_9 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h4;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] icmp_exitcond14549: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_6(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_8;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_9;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_10;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_12;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_13;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_14;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_50: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_50: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg [4:0] in_data_R_1_taskID; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_2;
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_3;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_4;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_5;
  reg [4:0] enable_R_taskID; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_6;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_7;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_8;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_9;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_10;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_11;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_12;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_17; // @[Bitwise.scala 108:18]
  wire  _T_18; // @[Bitwise.scala 108:44]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [4:0] task_input; // @[PhiNode.scala 250:43]
  wire [4:0] _GEN_18; // @[PhiNode.scala 253:20]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_13;
  wire  _T_22; // @[Conditional.scala 37:30]
  wire  _T_23; // @[PhiNode.scala 268:37]
  wire  _T_24; // @[PhiNode.scala 277:27]
  wire  _T_25; // @[PhiNode.scala 283:19]
  wire  _T_26; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_30; // @[PhiNode.scala 283:19]
  wire  _GEN_33; // @[PhiNode.scala 277:46]
  wire  _T_29; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_58; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_60; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_91; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_93; // @[Conditional.scala 39:67]
  wire  _GEN_113; // @[PhiNode.scala 283:19]
  wire  _GEN_114; // @[PhiNode.scala 283:19]
  wire  _GEN_116; // @[PhiNode.scala 291:19]
  wire  _GEN_117; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_17 = mask_R[0]; // @[Bitwise.scala 108:18]
  assign _T_18 = mask_R[1]; // @[Bitwise.scala 108:44]
  assign _T_19 = {_T_17,_T_18}; // @[Cat.scala 29:58]
  assign sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[PhiNode.scala 250:43]
  assign _GEN_18 = sel ? in_data_R_1_taskID : in_data_R_0_taskID; // @[PhiNode.scala 253:20]
  assign _GEN_19 = sel ? in_data_R_1_data : 32'h0; // @[PhiNode.scala 253:20]
  assign _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_20 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 265:74]
  assign _T_22 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_23 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_24 = enable_valid_R & _T_23; // @[PhiNode.scala 277:27]
  assign _T_25 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_26 = _T_25 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_30 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_33 = _T_24 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _T_29 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_58 = _T_33 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_60 = _T_33 ? task_input : _GEN_18; // @[Conditional.scala 39:67]
  assign _GEN_91 = _T_29 ? _GEN_19 : _GEN_58; // @[Conditional.scala 39:67]
  assign _GEN_93 = _T_29 ? _GEN_18 : _GEN_60; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_taskID = _T_22 ? _GEN_18 : _GEN_93; // @[PhiNode.scala 253:20 PhiNode.scala 327:44]
  assign io_Out_0_bits_data = _T_22 ? _GEN_19 : _GEN_91; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_113 = _T_22 & _T_24; // @[PhiNode.scala 283:19]
  assign _GEN_114 = _GEN_113 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_116 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_117 = _GEN_113 & _GEN_116; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_taskID = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  enable_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  enable_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mask_R = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mask_valid_R = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fire_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  state = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_22) begin
        if (_T_14) begin
          in_data_R_0_taskID <= io_InData_0_bits_taskID;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_14) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              in_data_R_0_taskID <= 5'h0;
            end else begin
              if (_T_14) begin
                in_data_R_0_taskID <= io_InData_0_bits_taskID;
              end
            end
          end else begin
            if (_T_14) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_taskID <= 5'h0;
    end else begin
      if (_T_22) begin
        if (_T_16) begin
          in_data_R_1_taskID <= io_InData_1_bits_taskID;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            in_data_R_1_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_taskID <= io_InData_1_bits_taskID;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              in_data_R_1_taskID <= 5'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_taskID <= io_InData_1_bits_taskID;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_taskID <= io_InData_1_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_22) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_22) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_22) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_22) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_12) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_22) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_22) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_22) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_22) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_22) begin
        out_valid_R_0 <= _GEN_33;
      end else begin
        if (_T_20) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_22) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_22) begin
        if (_T_24) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_dw_conv_013551: Output fired @ %d, Value: %d\n",_GEN_30,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_117 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_dw_conv_013551: Output flushed @ %d, Value: %d\n",_GEN_30,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_6(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_4;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_5;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_6;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_7;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_8;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_9;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_10;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_11;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_17; // @[Bitwise.scala 108:18]
  wire  _T_18; // @[Bitwise.scala 108:44]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_12;
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _T_25; // @[PhiNode.scala 268:37]
  wire  _T_26; // @[PhiNode.scala 277:27]
  wire  _T_27; // @[PhiNode.scala 283:19]
  wire  _T_28; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_32; // @[PhiNode.scala 283:19]
  wire  _GEN_35; // @[PhiNode.scala 277:46]
  wire  _GEN_36; // @[PhiNode.scala 277:46]
  wire  _T_31; // @[Conditional.scala 37:30]
  wire  _T_32; // @[PhiNode.scala 299:31]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_70; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_108; // @[Conditional.scala 39:67]
  wire  _GEN_138; // @[PhiNode.scala 283:19]
  wire  _GEN_139; // @[PhiNode.scala 283:19]
  wire  _GEN_141; // @[PhiNode.scala 291:19]
  wire  _GEN_142; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_17 = mask_R[0]; // @[Bitwise.scala 108:18]
  assign _T_18 = mask_R[1]; // @[Bitwise.scala 108:44]
  assign _T_19 = {_T_17,_T_18}; // @[Cat.scala 29:58]
  assign sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  assign _GEN_19 = sel ? in_data_R_1_data : 32'h0; // @[PhiNode.scala 253:20]
  assign _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_20 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = _T_21 | fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 265:74]
  assign _T_24 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_25 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_26 = enable_valid_R & _T_25; // @[PhiNode.scala 277:27]
  assign _T_27 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_28 = _T_27 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_32 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_35 = _T_26 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_36 = _T_26 | _GEN_23; // @[PhiNode.scala 277:46]
  assign _T_31 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_32 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_70 = _T_36 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_108 = _T_31 ? _GEN_19 : _GEN_70; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_24 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_data = _T_24 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_138 = _T_24 & _T_26; // @[PhiNode.scala 283:19]
  assign _GEN_139 = _GEN_138 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_141 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_142 = _GEN_138 & _GEN_141; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mask_R = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mask_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fire_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  fire_R_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_24) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_24) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_0 <= _GEN_35;
      end else begin
        if (_T_20) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_1 <= _GEN_36;
      end else begin
        if (_T_21) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        fire_R_1 <= _GEN_22;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            fire_R_1 <= 1'h0;
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_1 <= 1'h0;
            end else begin
              fire_R_1 <= _GEN_22;
            end
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_139 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_dw_conv_s1_r_dw__y_013452: Output fired @ %d, Value: %d\n",_GEN_32,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_142 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_dw_conv_s1_r_dw__y_013452: Output flushed @ %d, Value: %d\n",_GEN_32,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_26(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add2853: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_27(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_7 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_mul2954: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_28(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add3055: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_8(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_56: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [UBR] br_56: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_7(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  input  [31:0] io_InData_0_bits_data,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [4:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg [31:0] in_data_R_0_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_6;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_7;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_8;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_9;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_10;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire [4:0] task_input; // @[PhiNode.scala 250:43]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_10; // @[PhiNode.scala 258:26]
  wire  _GEN_11; // @[PhiNode.scala 258:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_12; // @[PhiNode.scala 258:26]
  wire  _GEN_13; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_11;
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[PhiNode.scala 277:27]
  wire  _T_20; // @[PhiNode.scala 283:19]
  wire  _T_21; // @[PhiNode.scala 283:19]
  wire  _GEN_15; // @[PhiNode.scala 277:46]
  wire  _GEN_16; // @[PhiNode.scala 277:46]
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _T_25; // @[PhiNode.scala 299:31]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_42; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_44; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_69; // @[Conditional.scala 39:67]
  wire [4:0] _GEN_71; // @[Conditional.scala 39:67]
  wire  _GEN_89; // @[PhiNode.scala 283:19]
  wire  _GEN_90; // @[PhiNode.scala 283:19]
  wire  _GEN_92; // @[PhiNode.scala 291:19]
  wire  _GEN_93; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_11 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_13 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_13 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[PhiNode.scala 250:43]
  assign _T_14 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_10 = _T_14 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_11 = _T_14 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_15 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_12 = _T_15 | fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_13 = _T_15 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_14; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_15; // @[PhiNode.scala 265:74]
  assign _T_18 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & in_data_valid_R_0; // @[PhiNode.scala 277:27]
  assign _T_20 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_21 = _T_20 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_15 = _T_19 | _GEN_11; // @[PhiNode.scala 277:46]
  assign _GEN_16 = _T_19 | _GEN_13; // @[PhiNode.scala 277:46]
  assign _T_24 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_25 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_28 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_42 = _T_28 ? 32'h0 : in_data_R_0_data; // @[Conditional.scala 39:67]
  assign _GEN_44 = _T_28 ? task_input : in_data_R_0_taskID; // @[Conditional.scala 39:67]
  assign _GEN_69 = _T_24 ? in_data_R_0_data : _GEN_42; // @[Conditional.scala 39:67]
  assign _GEN_71 = _T_24 ? in_data_R_0_taskID : _GEN_44; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_taskID = _T_18 ? in_data_R_0_taskID : _GEN_71; // @[PhiNode.scala 253:20 PhiNode.scala 327:44]
  assign io_Out_0_bits_data = _T_18 ? in_data_R_0_data : _GEN_69; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_taskID = _T_18 ? in_data_R_0_taskID : _GEN_71; // @[PhiNode.scala 253:20 PhiNode.scala 327:44]
  assign io_Out_1_bits_data = _T_18 ? in_data_R_0_data : _GEN_69; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_89 = _T_18 & _T_19; // @[PhiNode.scala 283:19]
  assign _GEN_90 = _GEN_89 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_92 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_93 = _GEN_89 & _GEN_92; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fire_R_1 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_18) begin
        if (_T_13) begin
          in_data_R_0_taskID <= io_InData_0_bits_taskID;
        end
      end else begin
        if (_T_24) begin
          if (_T_25) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_13) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end else begin
          if (_T_28) begin
            if (_T_25) begin
              in_data_R_0_taskID <= 5'h0;
            end else begin
              if (_T_13) begin
                in_data_R_0_taskID <= io_InData_0_bits_taskID;
              end
            end
          end else begin
            if (_T_13) begin
              in_data_R_0_taskID <= io_InData_0_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_data <= 32'h0;
    end else begin
      if (_T_18) begin
        if (_T_13) begin
          in_data_R_0_data <= io_InData_0_bits_data;
        end
      end else begin
        if (_T_24) begin
          if (_T_25) begin
            in_data_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end else begin
          if (_T_28) begin
            if (_T_25) begin
              in_data_R_0_data <= 32'h0;
            end else begin
              if (_T_13) begin
                in_data_R_0_data <= io_InData_0_bits_data;
              end
            end
          end else begin
            if (_T_13) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_24) begin
          if (_T_25) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_28) begin
            if (_T_25) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_18) begin
        if (_T_11) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_24) begin
          if (_T_25) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_28) begin
            if (_T_25) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_11) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_11) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_11) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_24) begin
          if (_T_25) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_11) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_28) begin
            if (_T_25) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_11) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_11) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_24) begin
          if (_T_25) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_28) begin
            if (_T_25) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        out_valid_R_0 <= _GEN_15;
      end else begin
        if (_T_14) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        out_valid_R_1 <= _GEN_16;
      end else begin
        if (_T_15) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        fire_R_0 <= _GEN_10;
      end else begin
        if (_T_24) begin
          if (_T_25) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_10;
          end
        end else begin
          if (_T_28) begin
            if (_T_25) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_10;
            end
          end else begin
            fire_R_0 <= _GEN_10;
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        fire_R_1 <= _GEN_12;
      end else begin
        if (_T_24) begin
          if (_T_25) begin
            fire_R_1 <= 1'h0;
          end else begin
            fire_R_1 <= _GEN_12;
          end
        end else begin
          if (_T_28) begin
            if (_T_25) begin
              fire_R_1 <= 1'h0;
            end else begin
              fire_R_1 <= _GEN_12;
            end
          end else begin
            fire_R_1 <= _GEN_12;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_18) begin
        if (_T_19) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_24) begin
          if (_T_25) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_28) begin
            if (_T_25) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_90 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phiadd38_lcssa57: Output fired @ %d, Value: %d\n",io_InData_0_bits_taskID,value,in_data_R_0_data); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_93 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phiadd38_lcssa57: Output flushed @ %d, Value: %d\n",io_InData_0_bits_taskID,value,in_data_R_0_data); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_29(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_inc4158: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_30(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_9 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h3;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] icmp_exitcond14459: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_7(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_8;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_9;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_10;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_12;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_13;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_14;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_60: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_60: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_8(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  input  [31:0] io_InData_0_bits_data,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_0_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_6;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_7;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_8;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_9;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_10;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_17; // @[Bitwise.scala 108:18]
  wire  _T_18; // @[Bitwise.scala 108:44]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_11;
  wire  _T_22; // @[Conditional.scala 37:30]
  wire  _T_23; // @[PhiNode.scala 268:37]
  wire  _T_24; // @[PhiNode.scala 277:27]
  wire  _T_25; // @[PhiNode.scala 283:19]
  wire  _T_26; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_30; // @[PhiNode.scala 283:19]
  wire  _GEN_33; // @[PhiNode.scala 277:46]
  wire  _T_29; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_58; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_91; // @[Conditional.scala 39:67]
  wire  _GEN_113; // @[PhiNode.scala 283:19]
  wire  _GEN_114; // @[PhiNode.scala 283:19]
  wire  _GEN_116; // @[PhiNode.scala 291:19]
  wire  _GEN_117; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_17 = mask_R[0]; // @[Bitwise.scala 108:18]
  assign _T_18 = mask_R[1]; // @[Bitwise.scala 108:44]
  assign _T_19 = {_T_17,_T_18}; // @[Cat.scala 29:58]
  assign sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  assign _GEN_19 = sel ? in_data_R_1_data : in_data_R_0_data; // @[PhiNode.scala 253:20]
  assign _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_20 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 265:74]
  assign _T_22 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_23 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_24 = enable_valid_R & _T_23; // @[PhiNode.scala 277:27]
  assign _T_25 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_26 = _T_25 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_30 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_33 = _T_24 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _T_29 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_58 = _T_33 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_91 = _T_29 ? _GEN_19 : _GEN_58; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_22 ? _GEN_19 : _GEN_91; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_113 = _T_22 & _T_24; // @[PhiNode.scala 283:19]
  assign _GEN_114 = _GEN_113 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_116 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_117 = _GEN_113 & _GEN_116; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mask_R = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mask_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fire_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_data <= 32'h0;
    end else begin
      if (_T_22) begin
        if (_T_14) begin
          in_data_R_0_data <= io_InData_0_bits_data;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            in_data_R_0_data <= 32'h0;
          end else begin
            if (_T_14) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              in_data_R_0_data <= 32'h0;
            end else begin
              if (_T_14) begin
                in_data_R_0_data <= io_InData_0_bits_data;
              end
            end
          end else begin
            if (_T_14) begin
              in_data_R_0_data <= io_InData_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_22) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_22) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_22) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_22) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_22) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_22) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_22) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_22) begin
        out_valid_R_0 <= _GEN_33;
      end else begin
        if (_T_20) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_22) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_22) begin
        if (_T_24) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_29) begin
          if (fire_mask_0) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_33) begin
            if (fire_mask_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_114 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_dw_conv_113361: Output fired @ %d, Value: %d\n",_GEN_30,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_117 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_dw_conv_113361: Output flushed @ %d, Value: %d\n",_GEN_30,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_9(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_4;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_5;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_6;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_7;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_8;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_9;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_10;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_11;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_17; // @[Bitwise.scala 108:18]
  wire  _T_18; // @[Bitwise.scala 108:44]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_12;
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _T_25; // @[PhiNode.scala 268:37]
  wire  _T_26; // @[PhiNode.scala 277:27]
  wire  _T_27; // @[PhiNode.scala 283:19]
  wire  _T_28; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_32; // @[PhiNode.scala 283:19]
  wire  _GEN_35; // @[PhiNode.scala 277:46]
  wire  _GEN_36; // @[PhiNode.scala 277:46]
  wire  _T_31; // @[Conditional.scala 37:30]
  wire  _T_32; // @[PhiNode.scala 299:31]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_70; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_108; // @[Conditional.scala 39:67]
  wire  _GEN_138; // @[PhiNode.scala 283:19]
  wire  _GEN_139; // @[PhiNode.scala 283:19]
  wire  _GEN_141; // @[PhiNode.scala 291:19]
  wire  _GEN_142; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_17 = mask_R[0]; // @[Bitwise.scala 108:18]
  assign _T_18 = mask_R[1]; // @[Bitwise.scala 108:44]
  assign _T_19 = {_T_17,_T_18}; // @[Cat.scala 29:58]
  assign sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  assign _GEN_19 = sel ? in_data_R_1_data : 32'h0; // @[PhiNode.scala 253:20]
  assign _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_20 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = _T_21 | fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 265:74]
  assign _T_24 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_25 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_26 = enable_valid_R & _T_25; // @[PhiNode.scala 277:27]
  assign _T_27 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_28 = _T_27 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_32 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_35 = _T_26 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_36 = _T_26 | _GEN_23; // @[PhiNode.scala 277:46]
  assign _T_31 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_32 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_70 = _T_36 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_108 = _T_31 ? _GEN_19 : _GEN_70; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_24 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_data = _T_24 ? _GEN_19 : _GEN_108; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_138 = _T_24 & _T_26; // @[PhiNode.scala 283:19]
  assign _GEN_139 = _GEN_138 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_141 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_142 = _GEN_138 & _GEN_141; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mask_R = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mask_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  fire_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  fire_R_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_24) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_24) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_0 <= _GEN_35;
      end else begin
        if (_T_20) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        out_valid_R_1 <= _GEN_36;
      end else begin
        if (_T_21) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        fire_R_1 <= _GEN_22;
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            fire_R_1 <= 1'h0;
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              fire_R_1 <= 1'h0;
            end else begin
              fire_R_1 <= _GEN_22;
            end
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_31) begin
          if (_T_32) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_36) begin
            if (_T_32) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_139 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_dw_conv_s1_r_dw__x_013262: Output fired @ %d, Value: %d\n",_GEN_32,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_142 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [PHI] phi_dw_conv_s1_r_dw__x_013262: Output flushed @ %d, Value: %d\n",_GEN_32,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_31(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add3563: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [GEP] Gep_arrayidx64: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOAD] ld_65: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOAD] ld_65: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [LOAD] ld_65: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SextNode_1(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[SextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[SextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[SextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[SextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[SextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[SextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[SextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[SextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[SextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[SextNode.scala 84:26]
  wire  _GEN_9; // @[SextNode.scala 84:26]
  wire  fire_mask_0; // @[SextNode.scala 90:74]
  reg  state; // @[SextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[SextNode.scala 93:27]
  wire  _T_16; // @[SextNode.scala 97:26]
  wire  _T_17; // @[SextNode.scala 110:28]
  wire  _T_18; // @[SextNode.scala 117:17]
  wire  _T_19; // @[SextNode.scala 117:17]
  wire  _GEN_10; // @[SextNode.scala 110:47]
  wire  _GEN_11; // @[SextNode.scala 110:47]
  wire  _GEN_42; // @[SextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[SextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[SextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[SextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[SextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[SextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[SextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[SextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[SextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[SextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[SextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[SextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[SextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[SextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[SextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[SextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[SextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[SextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[SextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] sextconv3766: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[SextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_32(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [4:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_add3867: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_33(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] binaryOp_inc68: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_34(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_9 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h3;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [COMPUTE] icmp_exitcond69: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_8(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_8;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_9;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_10;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_12;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_13;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_14;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_70: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CBR] br_70: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const0: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_1(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const1: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_2(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const2: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_3(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [4:0] io_Out_bits_taskID
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign io_Out_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 126:15]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const3: Output fired @ %d, Value: %d\n",taskID,value,32'sh0); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_4(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const4: Output fired @ %d, Value: %d\n",taskID,value,32'sh3); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_5(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const5: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_6(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const6: Output fired @ %d, Value: %d\n",taskID,value,32'sh4); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_7(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [4:0] io_Out_bits_taskID
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign io_Out_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 126:15]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const7: Output fired @ %d, Value: %d\n",taskID,value,32'sh0); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_8(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [4:0] io_Out_bits_taskID
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign io_Out_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 126:15]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const8: Output fired @ %d, Value: %d\n",taskID,value,32'sh0); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_9(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const9: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_10(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const10: Output fired @ %d, Value: %d\n",taskID,value,32'sh3); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_11(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [4:0] io_Out_bits_taskID
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign io_Out_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 126:15]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const11: Output fired @ %d, Value: %d\n",taskID,value,32'sh0); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_12(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const12: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_13(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_reduction] [TID->%d] [CONST] const13: Output fired @ %d, Value: %d\n",taskID,value,32'sh3); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module extracted_function_reductionDF(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [4:0]  io_in_bits_enable_taskID,
  input         io_in_bits_enable_control,
  input         io_in_bits_data_field10_predicate,
  input  [4:0]  io_in_bits_data_field10_taskID,
  input  [31:0] io_in_bits_data_field10_data,
  input         io_in_bits_data_field9_predicate,
  input  [4:0]  io_in_bits_data_field9_taskID,
  input  [31:0] io_in_bits_data_field9_data,
  input         io_in_bits_data_field8_predicate,
  input  [4:0]  io_in_bits_data_field8_taskID,
  input  [31:0] io_in_bits_data_field8_data,
  input         io_in_bits_data_field7_predicate,
  input  [4:0]  io_in_bits_data_field7_taskID,
  input  [31:0] io_in_bits_data_field7_data,
  input         io_in_bits_data_field6_predicate,
  input  [4:0]  io_in_bits_data_field6_taskID,
  input  [31:0] io_in_bits_data_field6_data,
  input         io_in_bits_data_field5_predicate,
  input  [4:0]  io_in_bits_data_field5_taskID,
  input  [31:0] io_in_bits_data_field5_data,
  input         io_in_bits_data_field4_predicate,
  input  [4:0]  io_in_bits_data_field4_taskID,
  input  [31:0] io_in_bits_data_field4_data,
  input         io_in_bits_data_field3_predicate,
  input  [4:0]  io_in_bits_data_field3_taskID,
  input  [31:0] io_in_bits_data_field3_data,
  input         io_in_bits_data_field2_predicate,
  input  [4:0]  io_in_bits_data_field2_taskID,
  input  [31:0] io_in_bits_data_field2_data,
  input         io_in_bits_data_field1_predicate,
  input  [4:0]  io_in_bits_data_field1_taskID,
  input  [31:0] io_in_bits_data_field1_data,
  input         io_in_bits_data_field0_predicate,
  input  [4:0]  io_in_bits_data_field0_taskID,
  input  [31:0] io_in_bits_data_field0_data,
  input         io_MemResp_valid,
  input         io_MemResp_bits_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemResp_bits_iswrite,
  input  [31:0] io_MemResp_bits_tile,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  output [31:0] io_MemReq_bits_tile,
  input         io_out_ready,
  output        io_out_valid,
  output [4:0]  io_out_bits_enable_taskID,
  output        io_out_bits_enable_control
);
  wire  MemCtrl_clock; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_reset; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_WriteIn_0_ready; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_WriteIn_0_valid; // @[extracted_function_reduction.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_0_bits_address; // @[extracted_function_reduction.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_0_bits_data; // @[extracted_function_reduction.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_0_bits_taskID; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_WriteOut_0_valid; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_ReadIn_0_ready; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_ReadIn_0_valid; // @[extracted_function_reduction.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_0_bits_address; // @[extracted_function_reduction.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_0_bits_taskID; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_ReadIn_1_ready; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_ReadIn_1_valid; // @[extracted_function_reduction.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_1_bits_address; // @[extracted_function_reduction.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_1_bits_taskID; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_ReadOut_0_valid; // @[extracted_function_reduction.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_0_data; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_ReadOut_1_valid; // @[extracted_function_reduction.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_1_data; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_MemResp_valid; // @[extracted_function_reduction.scala 45:23]
  wire [31:0] MemCtrl_io_MemResp_bits_data; // @[extracted_function_reduction.scala 45:23]
  wire [7:0] MemCtrl_io_MemResp_bits_tag; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_MemResp_bits_iswrite; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_MemReq_ready; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_MemReq_valid; // @[extracted_function_reduction.scala 45:23]
  wire [31:0] MemCtrl_io_MemReq_bits_addr; // @[extracted_function_reduction.scala 45:23]
  wire [31:0] MemCtrl_io_MemReq_bits_data; // @[extracted_function_reduction.scala 45:23]
  wire [3:0] MemCtrl_io_MemReq_bits_mask; // @[extracted_function_reduction.scala 45:23]
  wire [7:0] MemCtrl_io_MemReq_bits_tag; // @[extracted_function_reduction.scala 45:23]
  wire [4:0] MemCtrl_io_MemReq_bits_taskID; // @[extracted_function_reduction.scala 45:23]
  wire  MemCtrl_io_MemReq_bits_iswrite; // @[extracted_function_reduction.scala 45:23]
  wire  InputSplitter_clock; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_reset; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_In_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_In_valid; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_enable_taskID; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_In_bits_enable_control; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field10_data; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field9_data; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_data_field8_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field8_data; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field7_data; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_data_field6_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field6_data; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field5_data; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_data_field4_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field4_data; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field3_data; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field2_data; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_data_field1_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field1_data; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_data_field0_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field0_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_enable_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_enable_valid; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_Out_enable_bits_taskID; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_enable_bits_control; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field10_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field10_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field10_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field9_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field9_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field9_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field8_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field8_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field8_0_bits_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field8_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field8_1_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field8_1_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field8_1_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field8_2_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field8_2_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field8_2_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field7_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field7_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field7_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field7_1_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field7_1_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field7_1_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field6_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field6_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field6_0_bits_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field6_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field6_1_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field6_1_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field6_1_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field6_2_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field6_2_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field6_2_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field5_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field5_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field5_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field5_1_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field5_1_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field5_1_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field4_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field4_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field4_0_bits_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field4_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field4_1_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field4_1_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field4_1_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field4_2_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field4_2_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field4_2_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field3_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field3_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field3_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field2_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field2_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field2_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_0_bits_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field0_0_ready; // @[extracted_function_reduction.scala 53:29]
  wire  InputSplitter_io_Out_data_field0_0_valid; // @[extracted_function_reduction.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field0_0_bits_taskID; // @[extracted_function_reduction.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field0_0_bits_data; // @[extracted_function_reduction.scala 53:29]
  wire  Loop_0_clock; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_reset; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_enable_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_enable_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_enable_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_enable_bits_control; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_InLiveIn_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_0_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_InLiveIn_1_valid; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_1_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_InLiveIn_2_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_2_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_2_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field2_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field2_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field1_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field0_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field0_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_activate_loop_start_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_activate_loop_back_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_loopBack_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_loopBack_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_loopBack_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_loopBack_0_bits_control; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_loopFinish_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_loopFinish_0_bits_control; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_CarryDepenIn_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_CarryDepenIn_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_CarryDepenIn_0_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_CarryDepenIn_1_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_CarryDepenIn_1_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_CarryDepenIn_1_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_CarryDepenIn_1_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_CarryDepenOut_field1_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_CarryDepenOut_field1_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_CarryDepenOut_field1_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_CarryDepenOut_field1_0_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_CarryDepenOut_field0_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_InLiveOut_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_InLiveOut_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_InLiveOut_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_InLiveOut_0_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_OutLiveOut_field0_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_OutLiveOut_field0_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveOut_field0_0_bits_data; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_loopExit_0_ready; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_loopExit_0_valid; // @[extracted_function_reduction.scala 62:22]
  wire [4:0] Loop_0_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_0_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 62:22]
  wire  Loop_1_clock; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_reset; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_enable_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_enable_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_enable_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_enable_bits_control; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveIn_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveIn_1_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_1_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_1_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveIn_2_valid; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_2_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveIn_3_valid; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_3_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field3_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field2_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field1_0_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_activate_loop_start_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_activate_loop_back_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_loopBack_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_loopBack_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_loopBack_0_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_loopBack_0_bits_control; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_loopFinish_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_loopFinish_0_bits_control; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_CarryDepenIn_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_CarryDepenIn_0_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_CarryDepenIn_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_CarryDepenIn_1_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_CarryDepenIn_1_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_CarryDepenIn_1_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_CarryDepenIn_1_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_CarryDepenOut_field1_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_CarryDepenOut_field1_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_CarryDepenOut_field1_0_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_CarryDepenOut_field1_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_CarryDepenOut_field0_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveOut_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_InLiveOut_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_InLiveOut_0_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_InLiveOut_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveOut_field0_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_OutLiveOut_field0_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveOut_field0_0_bits_data; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_loopExit_0_ready; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_loopExit_0_valid; // @[extracted_function_reduction.scala 64:22]
  wire [4:0] Loop_1_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_1_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 64:22]
  wire  Loop_2_clock; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_reset; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_enable_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_enable_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_enable_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_enable_bits_control; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_0_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_1_valid; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_1_bits_predicate; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_InLiveIn_1_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_1_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_2_valid; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_2_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_3_valid; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_3_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_4_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_4_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_InLiveIn_4_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_4_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_5_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_InLiveIn_5_valid; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_InLiveIn_5_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field5_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field5_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field4_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field4_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field3_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field2_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field1_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field1_0_bits_predicate; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_OutLiveIn_field1_0_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field1_1_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field1_1_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_OutLiveIn_field1_1_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field1_1_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field0_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_activate_loop_start_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_activate_loop_back_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_loopBack_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_loopBack_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_loopBack_0_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_loopBack_0_bits_control; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_loopFinish_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_loopFinish_0_bits_control; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_CarryDepenIn_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_CarryDepenIn_0_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_CarryDepenIn_0_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_CarryDepenOut_field0_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire [31:0] Loop_2_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_loopExit_0_ready; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_loopExit_0_valid; // @[extracted_function_reduction.scala 66:22]
  wire [4:0] Loop_2_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_2_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 66:22]
  wire  Loop_3_clock; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_reset; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_enable_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_enable_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_enable_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_enable_bits_control; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_1_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_1_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_2_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_2_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_3_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_3_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_4_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_4_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_InLiveIn_4_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_4_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_5_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_5_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_InLiveIn_5_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_5_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_6_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_6_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_6_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_7_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_7_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_7_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_8_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_InLiveIn_8_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_InLiveIn_8_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_InLiveIn_8_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field8_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field8_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field8_1_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field8_1_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field8_1_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field7_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field7_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field6_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field6_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field5_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field5_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_OutLiveIn_field5_0_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field4_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field4_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field3_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field2_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field1_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field0_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_activate_loop_start_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_activate_loop_back_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_loopBack_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_loopBack_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_loopBack_0_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_loopBack_0_bits_control; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_loopFinish_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_loopFinish_0_bits_control; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_CarryDepenIn_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_CarryDepenIn_0_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_CarryDepenIn_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_CarryDepenOut_field0_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire [31:0] Loop_3_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_loopExit_0_ready; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_loopExit_0_valid; // @[extracted_function_reduction.scala 68:22]
  wire [4:0] Loop_3_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_3_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 68:22]
  wire  Loop_4_clock; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_reset; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_enable_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_enable_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_enable_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_enable_bits_control; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_1_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_1_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_2_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_2_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_3_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_InLiveIn_3_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_3_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_4_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_4_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_InLiveIn_4_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_4_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_5_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_5_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_5_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_6_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_6_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_6_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_7_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_7_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_InLiveIn_7_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_7_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_8_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_8_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_InLiveIn_8_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_8_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_9_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_9_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_9_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_10_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_10_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_InLiveIn_10_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_10_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_11_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_InLiveIn_11_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_InLiveIn_11_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field11_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field11_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field11_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field10_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field10_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_OutLiveIn_field10_0_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field10_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field10_1_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field10_1_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field10_1_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field9_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field9_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field9_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field8_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field8_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field7_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field7_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_OutLiveIn_field7_0_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field6_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field6_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field5_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field5_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field4_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field4_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field3_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_OutLiveIn_field3_0_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field2_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field1_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field0_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_activate_loop_start_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_activate_loop_back_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_loopBack_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_loopBack_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_loopBack_0_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_loopBack_0_bits_control; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_loopFinish_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_loopFinish_0_bits_control; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_CarryDepenIn_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_CarryDepenIn_0_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_CarryDepenIn_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_CarryDepenOut_field0_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire [31:0] Loop_4_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_loopExit_0_ready; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_loopExit_0_valid; // @[extracted_function_reduction.scala 70:22]
  wire [4:0] Loop_4_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_4_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 70:22]
  wire  Loop_5_clock; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_reset; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_enable_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_enable_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_enable_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_enable_bits_control; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_InLiveIn_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_1_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_1_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_2_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_InLiveIn_2_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_2_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_3_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_InLiveIn_3_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_3_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_4_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_4_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_InLiveIn_4_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_4_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_5_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_5_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_5_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_6_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_6_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_InLiveIn_6_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_6_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_7_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_7_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_7_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_8_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_8_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_InLiveIn_8_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_8_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_9_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_9_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_9_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_10_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_10_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_10_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_11_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_11_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_InLiveIn_11_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_11_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_12_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_12_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_12_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_13_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_13_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_13_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_14_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_InLiveIn_14_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_InLiveIn_14_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field14_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field14_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field14_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field13_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field13_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field13_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field12_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field12_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field12_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field11_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field11_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_OutLiveIn_field11_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field11_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field10_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field10_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field10_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field9_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field9_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field9_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field8_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field8_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field7_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field7_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field6_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field6_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_OutLiveIn_field6_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field5_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field5_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field4_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field4_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field3_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_OutLiveIn_field3_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field2_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_OutLiveIn_field2_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field1_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field0_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_OutLiveIn_field0_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field0_1_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_OutLiveIn_field0_1_valid; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_OutLiveIn_field0_1_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_activate_loop_start_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_activate_loop_back_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_loopBack_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_loopBack_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_loopBack_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_loopBack_0_bits_control; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_loopFinish_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_loopFinish_0_bits_control; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_CarryDepenIn_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_CarryDepenIn_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_CarryDepenIn_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_CarryDepenOut_field0_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire [31:0] Loop_5_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_loopExit_0_ready; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_loopExit_0_valid; // @[extracted_function_reduction.scala 72:22]
  wire [4:0] Loop_5_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 72:22]
  wire  Loop_5_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 72:22]
  wire  bb_entry0_clock; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_reset; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 80:25]
  wire [4:0] bb_entry0_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_Out_0_ready; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_Out_0_valid; // @[extracted_function_reduction.scala 80:25]
  wire [4:0] bb_entry0_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_Out_0_bits_control; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_Out_1_ready; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_Out_1_valid; // @[extracted_function_reduction.scala 80:25]
  wire [4:0] bb_entry0_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_Out_1_bits_control; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_Out_2_ready; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_Out_2_valid; // @[extracted_function_reduction.scala 80:25]
  wire [4:0] bb_entry0_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 80:25]
  wire  bb_entry0_io_Out_2_bits_control; // @[extracted_function_reduction.scala 80:25]
  wire  bb_for_body_lr_ph1_clock; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_reset; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 82:34]
  wire [4:0] bb_for_body_lr_ph1_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_0_ready; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_0_valid; // @[extracted_function_reduction.scala 82:34]
  wire [4:0] bb_for_body_lr_ph1_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_0_bits_control; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_1_ready; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_1_valid; // @[extracted_function_reduction.scala 82:34]
  wire [4:0] bb_for_body_lr_ph1_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_1_bits_control; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_2_ready; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_2_valid; // @[extracted_function_reduction.scala 82:34]
  wire [4:0] bb_for_body_lr_ph1_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_2_bits_control; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_3_ready; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_3_valid; // @[extracted_function_reduction.scala 82:34]
  wire [4:0] bb_for_body_lr_ph1_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_3_bits_control; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_4_ready; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_4_valid; // @[extracted_function_reduction.scala 82:34]
  wire [4:0] bb_for_body_lr_ph1_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_body_lr_ph1_io_Out_4_bits_control; // @[extracted_function_reduction.scala 82:34]
  wire  bb_for_cond_cleanup_loopexit2_clock; // @[extracted_function_reduction.scala 84:45]
  wire  bb_for_cond_cleanup_loopexit2_reset; // @[extracted_function_reduction.scala 84:45]
  wire  bb_for_cond_cleanup_loopexit2_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 84:45]
  wire  bb_for_cond_cleanup_loopexit2_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 84:45]
  wire [4:0] bb_for_cond_cleanup_loopexit2_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 84:45]
  wire  bb_for_cond_cleanup_loopexit2_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 84:45]
  wire  bb_for_cond_cleanup_loopexit2_io_Out_0_ready; // @[extracted_function_reduction.scala 84:45]
  wire  bb_for_cond_cleanup_loopexit2_io_Out_0_valid; // @[extracted_function_reduction.scala 84:45]
  wire [4:0] bb_for_cond_cleanup_loopexit2_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 84:45]
  wire  bb_for_cond_cleanup_loopexit2_io_Out_0_bits_control; // @[extracted_function_reduction.scala 84:45]
  wire  bb_for_cond_cleanup3_clock; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_reset; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 86:36]
  wire [4:0] bb_for_cond_cleanup3_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_io_predicateIn_1_valid; // @[extracted_function_reduction.scala 86:36]
  wire [4:0] bb_for_cond_cleanup3_io_predicateIn_1_bits_taskID; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_io_predicateIn_1_bits_control; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_io_Out_0_ready; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_io_Out_0_valid; // @[extracted_function_reduction.scala 86:36]
  wire [4:0] bb_for_cond_cleanup3_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_cond_cleanup3_io_Out_0_bits_control; // @[extracted_function_reduction.scala 86:36]
  wire  bb_for_body4_clock; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_reset; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_MaskBB_0_ready; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 88:28]
  wire [1:0] bb_for_body4_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_0_ready; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_0_valid; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_0_bits_control; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_1_ready; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_1_valid; // @[extracted_function_reduction.scala 88:28]
  wire [4:0] bb_for_body4_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_1_bits_control; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_2_ready; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_2_valid; // @[extracted_function_reduction.scala 88:28]
  wire [4:0] bb_for_body4_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_2_bits_control; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_3_ready; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_3_valid; // @[extracted_function_reduction.scala 88:28]
  wire [4:0] bb_for_body4_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_Out_3_bits_control; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 88:28]
  wire [4:0] bb_for_body4_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_predicateIn_1_valid; // @[extracted_function_reduction.scala 88:28]
  wire [4:0] bb_for_body4_io_predicateIn_1_bits_taskID; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body4_io_predicateIn_1_bits_control; // @[extracted_function_reduction.scala 88:28]
  wire  bb_for_body7_preheader5_clock; // @[extracted_function_reduction.scala 90:39]
  wire  bb_for_body7_preheader5_reset; // @[extracted_function_reduction.scala 90:39]
  wire  bb_for_body7_preheader5_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 90:39]
  wire  bb_for_body7_preheader5_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 90:39]
  wire [4:0] bb_for_body7_preheader5_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 90:39]
  wire  bb_for_body7_preheader5_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 90:39]
  wire  bb_for_body7_preheader5_io_Out_0_ready; // @[extracted_function_reduction.scala 90:39]
  wire  bb_for_body7_preheader5_io_Out_0_valid; // @[extracted_function_reduction.scala 90:39]
  wire [4:0] bb_for_body7_preheader5_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 90:39]
  wire  bb_for_body7_preheader5_io_Out_0_bits_control; // @[extracted_function_reduction.scala 90:39]
  wire  bb_for_cond_cleanup6_loopexit6_clock; // @[extracted_function_reduction.scala 92:46]
  wire  bb_for_cond_cleanup6_loopexit6_reset; // @[extracted_function_reduction.scala 92:46]
  wire  bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 92:46]
  wire  bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 92:46]
  wire [4:0] bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 92:46]
  wire  bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 92:46]
  wire  bb_for_cond_cleanup6_loopexit6_io_Out_0_ready; // @[extracted_function_reduction.scala 92:46]
  wire  bb_for_cond_cleanup6_loopexit6_io_Out_0_valid; // @[extracted_function_reduction.scala 92:46]
  wire [4:0] bb_for_cond_cleanup6_loopexit6_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 92:46]
  wire  bb_for_cond_cleanup6_loopexit6_io_Out_0_bits_control; // @[extracted_function_reduction.scala 92:46]
  wire  bb_for_cond_cleanup67_clock; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_reset; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 94:37]
  wire [4:0] bb_for_cond_cleanup67_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_predicateIn_1_valid; // @[extracted_function_reduction.scala 94:37]
  wire [4:0] bb_for_cond_cleanup67_io_predicateIn_1_bits_taskID; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_predicateIn_1_bits_control; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_0_ready; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_0_valid; // @[extracted_function_reduction.scala 94:37]
  wire [4:0] bb_for_cond_cleanup67_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_1_ready; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_1_valid; // @[extracted_function_reduction.scala 94:37]
  wire [4:0] bb_for_cond_cleanup67_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_1_bits_control; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_2_ready; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_2_valid; // @[extracted_function_reduction.scala 94:37]
  wire [4:0] bb_for_cond_cleanup67_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_2_bits_control; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_3_ready; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_3_valid; // @[extracted_function_reduction.scala 94:37]
  wire [4:0] bb_for_cond_cleanup67_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_cond_cleanup67_io_Out_3_bits_control; // @[extracted_function_reduction.scala 94:37]
  wire  bb_for_body78_clock; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_reset; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_MaskBB_0_ready; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 96:29]
  wire [1:0] bb_for_body78_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_Out_0_ready; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_Out_0_valid; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_Out_0_bits_control; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_Out_1_ready; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_Out_1_valid; // @[extracted_function_reduction.scala 96:29]
  wire [4:0] bb_for_body78_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_Out_1_bits_control; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 96:29]
  wire [4:0] bb_for_body78_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_predicateIn_1_valid; // @[extracted_function_reduction.scala 96:29]
  wire [4:0] bb_for_body78_io_predicateIn_1_bits_taskID; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body78_io_predicateIn_1_bits_control; // @[extracted_function_reduction.scala 96:29]
  wire  bb_for_body15_lr_ph9_clock; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_reset; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 98:36]
  wire [4:0] bb_for_body15_lr_ph9_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_0_ready; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_0_valid; // @[extracted_function_reduction.scala 98:36]
  wire [4:0] bb_for_body15_lr_ph9_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_0_bits_control; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_1_ready; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_1_valid; // @[extracted_function_reduction.scala 98:36]
  wire [4:0] bb_for_body15_lr_ph9_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_1_bits_control; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_2_ready; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_2_valid; // @[extracted_function_reduction.scala 98:36]
  wire [4:0] bb_for_body15_lr_ph9_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_2_bits_control; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_3_ready; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_3_valid; // @[extracted_function_reduction.scala 98:36]
  wire [4:0] bb_for_body15_lr_ph9_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_body15_lr_ph9_io_Out_3_bits_control; // @[extracted_function_reduction.scala 98:36]
  wire  bb_for_cond_cleanup14_loopexit10_clock; // @[extracted_function_reduction.scala 100:48]
  wire  bb_for_cond_cleanup14_loopexit10_reset; // @[extracted_function_reduction.scala 100:48]
  wire  bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 100:48]
  wire  bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 100:48]
  wire [4:0] bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 100:48]
  wire  bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 100:48]
  wire  bb_for_cond_cleanup14_loopexit10_io_Out_0_ready; // @[extracted_function_reduction.scala 100:48]
  wire  bb_for_cond_cleanup14_loopexit10_io_Out_0_valid; // @[extracted_function_reduction.scala 100:48]
  wire [4:0] bb_for_cond_cleanup14_loopexit10_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 100:48]
  wire  bb_for_cond_cleanup14_loopexit10_io_Out_0_bits_control; // @[extracted_function_reduction.scala 100:48]
  wire  bb_for_cond_cleanup1411_clock; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_reset; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 102:39]
  wire [4:0] bb_for_cond_cleanup1411_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_predicateIn_1_valid; // @[extracted_function_reduction.scala 102:39]
  wire [4:0] bb_for_cond_cleanup1411_io_predicateIn_1_bits_taskID; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_predicateIn_1_bits_control; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_0_ready; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_0_valid; // @[extracted_function_reduction.scala 102:39]
  wire [4:0] bb_for_cond_cleanup1411_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_1_ready; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_1_valid; // @[extracted_function_reduction.scala 102:39]
  wire [4:0] bb_for_cond_cleanup1411_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_1_bits_control; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_2_ready; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_2_valid; // @[extracted_function_reduction.scala 102:39]
  wire [4:0] bb_for_cond_cleanup1411_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_2_bits_control; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_3_ready; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_3_valid; // @[extracted_function_reduction.scala 102:39]
  wire [4:0] bb_for_cond_cleanup1411_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_cond_cleanup1411_io_Out_3_bits_control; // @[extracted_function_reduction.scala 102:39]
  wire  bb_for_body1512_clock; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_reset; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_MaskBB_0_ready; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 104:31]
  wire [1:0] bb_for_body1512_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_0_ready; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_0_valid; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_0_bits_control; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_1_ready; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_1_valid; // @[extracted_function_reduction.scala 104:31]
  wire [4:0] bb_for_body1512_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_1_bits_control; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_2_ready; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_2_valid; // @[extracted_function_reduction.scala 104:31]
  wire [4:0] bb_for_body1512_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_2_bits_control; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_3_ready; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_3_valid; // @[extracted_function_reduction.scala 104:31]
  wire [4:0] bb_for_body1512_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_3_bits_control; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_4_ready; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_4_valid; // @[extracted_function_reduction.scala 104:31]
  wire [4:0] bb_for_body1512_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_4_bits_control; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_5_ready; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_5_valid; // @[extracted_function_reduction.scala 104:31]
  wire [4:0] bb_for_body1512_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_Out_5_bits_control; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 104:31]
  wire [4:0] bb_for_body1512_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_predicateIn_1_valid; // @[extracted_function_reduction.scala 104:31]
  wire [4:0] bb_for_body1512_io_predicateIn_1_bits_taskID; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_body1512_io_predicateIn_1_bits_control; // @[extracted_function_reduction.scala 104:31]
  wire  bb_for_cond_cleanup2013_clock; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_reset; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 106:39]
  wire [4:0] bb_for_cond_cleanup2013_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_0_ready; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_0_valid; // @[extracted_function_reduction.scala 106:39]
  wire [4:0] bb_for_cond_cleanup2013_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_1_ready; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_1_valid; // @[extracted_function_reduction.scala 106:39]
  wire [4:0] bb_for_cond_cleanup2013_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_1_bits_control; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_2_ready; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_2_valid; // @[extracted_function_reduction.scala 106:39]
  wire [4:0] bb_for_cond_cleanup2013_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_2_bits_control; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_3_ready; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_3_valid; // @[extracted_function_reduction.scala 106:39]
  wire [4:0] bb_for_cond_cleanup2013_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_cond_cleanup2013_io_Out_3_bits_control; // @[extracted_function_reduction.scala 106:39]
  wire  bb_for_body2114_clock; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_reset; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_MaskBB_0_ready; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 108:31]
  wire [1:0] bb_for_body2114_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_0_ready; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_0_valid; // @[extracted_function_reduction.scala 108:31]
  wire [4:0] bb_for_body2114_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_1_ready; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_1_valid; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_1_bits_control; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_2_ready; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_2_valid; // @[extracted_function_reduction.scala 108:31]
  wire [4:0] bb_for_body2114_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_2_bits_control; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_3_ready; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_3_valid; // @[extracted_function_reduction.scala 108:31]
  wire [4:0] bb_for_body2114_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_3_bits_control; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_4_ready; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_4_valid; // @[extracted_function_reduction.scala 108:31]
  wire [4:0] bb_for_body2114_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_Out_4_bits_control; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 108:31]
  wire [4:0] bb_for_body2114_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_predicateIn_1_valid; // @[extracted_function_reduction.scala 108:31]
  wire [4:0] bb_for_body2114_io_predicateIn_1_bits_taskID; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_body2114_io_predicateIn_1_bits_control; // @[extracted_function_reduction.scala 108:31]
  wire  bb_for_cond_cleanup2615_clock; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_reset; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_0_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_0_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_1_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_1_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_2_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_2_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_3_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_3_valid; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_3_bits_control; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_4_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_4_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_4_bits_control; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_5_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_5_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_6_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_6_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_6_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_6_bits_control; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_7_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_7_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_7_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_7_bits_control; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_8_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_8_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_8_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_8_bits_control; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_9_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_9_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_9_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_9_bits_control; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_10_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_10_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_10_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_10_bits_control; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_11_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_11_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_Out_11_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_Out_11_bits_control; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 110:39]
  wire [4:0] bb_for_cond_cleanup2615_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_cond_cleanup2615_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 110:39]
  wire  bb_for_body2716_clock; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_reset; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_MaskBB_0_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 112:31]
  wire [1:0] bb_for_body2716_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_MaskBB_1_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_MaskBB_1_valid; // @[extracted_function_reduction.scala 112:31]
  wire [1:0] bb_for_body2716_io_MaskBB_1_bits; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_0_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_0_valid; // @[extracted_function_reduction.scala 112:31]
  wire [4:0] bb_for_body2716_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_1_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_1_valid; // @[extracted_function_reduction.scala 112:31]
  wire [4:0] bb_for_body2716_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_2_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_2_valid; // @[extracted_function_reduction.scala 112:31]
  wire [4:0] bb_for_body2716_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_2_bits_control; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_3_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_3_valid; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_3_bits_control; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_4_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_4_valid; // @[extracted_function_reduction.scala 112:31]
  wire [4:0] bb_for_body2716_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_4_bits_control; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_5_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_5_valid; // @[extracted_function_reduction.scala 112:31]
  wire [4:0] bb_for_body2716_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_5_bits_control; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_6_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_6_valid; // @[extracted_function_reduction.scala 112:31]
  wire [4:0] bb_for_body2716_io_Out_6_bits_taskID; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_6_bits_control; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_7_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_7_valid; // @[extracted_function_reduction.scala 112:31]
  wire [4:0] bb_for_body2716_io_Out_7_bits_taskID; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_Out_7_bits_control; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 112:31]
  wire [4:0] bb_for_body2716_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_predicateIn_1_valid; // @[extracted_function_reduction.scala 112:31]
  wire [4:0] bb_for_body2716_io_predicateIn_1_bits_taskID; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_body2716_io_predicateIn_1_bits_control; // @[extracted_function_reduction.scala 112:31]
  wire  bb_for_cond_cleanup3317_clock; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_reset; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_0_ready; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_0_valid; // @[extracted_function_reduction.scala 114:39]
  wire [4:0] bb_for_cond_cleanup3317_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_1_ready; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_1_valid; // @[extracted_function_reduction.scala 114:39]
  wire [4:0] bb_for_cond_cleanup3317_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_2_ready; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_2_valid; // @[extracted_function_reduction.scala 114:39]
  wire [4:0] bb_for_cond_cleanup3317_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_2_bits_control; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_3_ready; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_3_valid; // @[extracted_function_reduction.scala 114:39]
  wire [4:0] bb_for_cond_cleanup3317_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_3_bits_control; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_4_ready; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_4_valid; // @[extracted_function_reduction.scala 114:39]
  wire [4:0] bb_for_cond_cleanup3317_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_4_bits_control; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_5_ready; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_5_valid; // @[extracted_function_reduction.scala 114:39]
  wire [4:0] bb_for_cond_cleanup3317_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_Out_5_bits_control; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 114:39]
  wire [4:0] bb_for_cond_cleanup3317_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_cond_cleanup3317_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 114:39]
  wire  bb_for_body3418_clock; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_reset; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_MaskBB_0_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 116:31]
  wire [1:0] bb_for_body3418_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_MaskBB_1_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_MaskBB_1_valid; // @[extracted_function_reduction.scala 116:31]
  wire [1:0] bb_for_body3418_io_MaskBB_1_bits; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_0_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_0_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_1_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_1_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_2_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_2_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_3_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_3_valid; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_3_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_4_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_4_valid; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_4_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_5_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_5_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_5_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_6_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_6_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_6_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_6_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_7_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_7_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_7_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_7_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_8_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_8_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_8_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_9_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_9_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_9_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_9_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_10_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_10_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_10_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_10_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_11_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_11_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_11_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_11_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_12_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_12_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_Out_12_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_Out_12_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_predicateIn_0_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_predicateIn_0_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_predicateIn_0_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_predicateIn_1_valid; // @[extracted_function_reduction.scala 116:31]
  wire [4:0] bb_for_body3418_io_predicateIn_1_bits_taskID; // @[extracted_function_reduction.scala 116:31]
  wire  bb_for_body3418_io_predicateIn_1_bits_control; // @[extracted_function_reduction.scala 116:31]
  wire  binaryOp_add0_clock; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_reset; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_enable_ready; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_enable_valid; // @[extracted_function_reduction.scala 125:29]
  wire [4:0] binaryOp_add0_io_enable_bits_taskID; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_enable_bits_control; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_Out_0_ready; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_Out_0_valid; // @[extracted_function_reduction.scala 125:29]
  wire [31:0] binaryOp_add0_io_Out_0_bits_data; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_Out_1_ready; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_Out_1_valid; // @[extracted_function_reduction.scala 125:29]
  wire [31:0] binaryOp_add0_io_Out_1_bits_data; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_LeftIO_ready; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_LeftIO_valid; // @[extracted_function_reduction.scala 125:29]
  wire [31:0] binaryOp_add0_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_RightIO_ready; // @[extracted_function_reduction.scala 125:29]
  wire  binaryOp_add0_io_RightIO_valid; // @[extracted_function_reduction.scala 125:29]
  wire [31:0] binaryOp_add0_io_RightIO_bits_data; // @[extracted_function_reduction.scala 125:29]
  wire  icmp_cmp1421_clock; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_reset; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_io_enable_ready; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_io_enable_valid; // @[extracted_function_reduction.scala 128:28]
  wire [4:0] icmp_cmp1421_io_enable_bits_taskID; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_io_enable_bits_control; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_io_Out_0_ready; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_io_Out_0_valid; // @[extracted_function_reduction.scala 128:28]
  wire [4:0] icmp_cmp1421_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 128:28]
  wire [31:0] icmp_cmp1421_io_Out_0_bits_data; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_io_LeftIO_ready; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_io_LeftIO_valid; // @[extracted_function_reduction.scala 128:28]
  wire [31:0] icmp_cmp1421_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_io_RightIO_ready; // @[extracted_function_reduction.scala 128:28]
  wire  icmp_cmp1421_io_RightIO_valid; // @[extracted_function_reduction.scala 128:28]
  wire [31:0] icmp_cmp1421_io_RightIO_bits_data; // @[extracted_function_reduction.scala 128:28]
  wire  br_2_clock; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_reset; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_enable_ready; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_enable_valid; // @[extracted_function_reduction.scala 131:20]
  wire [4:0] br_2_io_enable_bits_taskID; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_enable_bits_control; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_CmpIO_ready; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_CmpIO_valid; // @[extracted_function_reduction.scala 131:20]
  wire [4:0] br_2_io_CmpIO_bits_taskID; // @[extracted_function_reduction.scala 131:20]
  wire [31:0] br_2_io_CmpIO_bits_data; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_TrueOutput_0_ready; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 131:20]
  wire [4:0] br_2_io_TrueOutput_0_bits_taskID; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_FalseOutput_0_ready; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 131:20]
  wire [4:0] br_2_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 131:20]
  wire  br_2_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 131:20]
  wire  binaryOp_add43_clock; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_reset; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_enable_ready; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_enable_valid; // @[extracted_function_reduction.scala 134:30]
  wire [4:0] binaryOp_add43_io_enable_bits_taskID; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_enable_bits_control; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_Out_0_ready; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_Out_0_valid; // @[extracted_function_reduction.scala 134:30]
  wire [31:0] binaryOp_add43_io_Out_0_bits_data; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_Out_1_ready; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_Out_1_valid; // @[extracted_function_reduction.scala 134:30]
  wire [31:0] binaryOp_add43_io_Out_1_bits_data; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_LeftIO_ready; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_LeftIO_valid; // @[extracted_function_reduction.scala 134:30]
  wire [31:0] binaryOp_add43_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_RightIO_ready; // @[extracted_function_reduction.scala 134:30]
  wire  binaryOp_add43_io_RightIO_valid; // @[extracted_function_reduction.scala 134:30]
  wire [31:0] binaryOp_add43_io_RightIO_bits_data; // @[extracted_function_reduction.scala 134:30]
  wire  icmp_cmp51394_clock; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_reset; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_io_enable_ready; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_io_enable_valid; // @[extracted_function_reduction.scala 137:29]
  wire [4:0] icmp_cmp51394_io_enable_bits_taskID; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_io_enable_bits_control; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_io_Out_0_ready; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_io_Out_0_valid; // @[extracted_function_reduction.scala 137:29]
  wire [4:0] icmp_cmp51394_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 137:29]
  wire [31:0] icmp_cmp51394_io_Out_0_bits_data; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_io_LeftIO_ready; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_io_LeftIO_valid; // @[extracted_function_reduction.scala 137:29]
  wire [31:0] icmp_cmp51394_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_io_RightIO_ready; // @[extracted_function_reduction.scala 137:29]
  wire  icmp_cmp51394_io_RightIO_valid; // @[extracted_function_reduction.scala 137:29]
  wire [31:0] icmp_cmp51394_io_RightIO_bits_data; // @[extracted_function_reduction.scala 137:29]
  wire  binaryOp_add125_clock; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_reset; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_enable_ready; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_enable_valid; // @[extracted_function_reduction.scala 140:31]
  wire [4:0] binaryOp_add125_io_enable_bits_taskID; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_enable_bits_control; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_Out_0_ready; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_Out_0_valid; // @[extracted_function_reduction.scala 140:31]
  wire [31:0] binaryOp_add125_io_Out_0_bits_data; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_Out_1_ready; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_Out_1_valid; // @[extracted_function_reduction.scala 140:31]
  wire [31:0] binaryOp_add125_io_Out_1_bits_data; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_LeftIO_ready; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_LeftIO_valid; // @[extracted_function_reduction.scala 140:31]
  wire [31:0] binaryOp_add125_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_RightIO_ready; // @[extracted_function_reduction.scala 140:31]
  wire  binaryOp_add125_io_RightIO_valid; // @[extracted_function_reduction.scala 140:31]
  wire [31:0] binaryOp_add125_io_RightIO_bits_data; // @[extracted_function_reduction.scala 140:31]
  wire  icmp_cmp131376_clock; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_reset; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_io_enable_ready; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_io_enable_valid; // @[extracted_function_reduction.scala 143:30]
  wire [4:0] icmp_cmp131376_io_enable_bits_taskID; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_io_enable_bits_control; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_io_Out_0_ready; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_io_Out_0_valid; // @[extracted_function_reduction.scala 143:30]
  wire [4:0] icmp_cmp131376_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 143:30]
  wire [31:0] icmp_cmp131376_io_Out_0_bits_data; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_io_LeftIO_ready; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_io_LeftIO_valid; // @[extracted_function_reduction.scala 143:30]
  wire [31:0] icmp_cmp131376_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_io_RightIO_ready; // @[extracted_function_reduction.scala 143:30]
  wire  icmp_cmp131376_io_RightIO_valid; // @[extracted_function_reduction.scala 143:30]
  wire [31:0] icmp_cmp131376_io_RightIO_bits_data; // @[extracted_function_reduction.scala 143:30]
  wire  br_7_clock; // @[extracted_function_reduction.scala 146:20]
  wire  br_7_reset; // @[extracted_function_reduction.scala 146:20]
  wire  br_7_io_enable_ready; // @[extracted_function_reduction.scala 146:20]
  wire  br_7_io_enable_valid; // @[extracted_function_reduction.scala 146:20]
  wire [4:0] br_7_io_enable_bits_taskID; // @[extracted_function_reduction.scala 146:20]
  wire  br_7_io_enable_bits_control; // @[extracted_function_reduction.scala 146:20]
  wire  br_7_io_Out_0_ready; // @[extracted_function_reduction.scala 146:20]
  wire  br_7_io_Out_0_valid; // @[extracted_function_reduction.scala 146:20]
  wire [4:0] br_7_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 146:20]
  wire  br_7_io_Out_0_bits_control; // @[extracted_function_reduction.scala 146:20]
  wire  br_8_clock; // @[extracted_function_reduction.scala 149:20]
  wire  br_8_reset; // @[extracted_function_reduction.scala 149:20]
  wire  br_8_io_enable_ready; // @[extracted_function_reduction.scala 149:20]
  wire  br_8_io_enable_valid; // @[extracted_function_reduction.scala 149:20]
  wire [4:0] br_8_io_enable_bits_taskID; // @[extracted_function_reduction.scala 149:20]
  wire  br_8_io_enable_bits_control; // @[extracted_function_reduction.scala 149:20]
  wire  br_8_io_Out_0_ready; // @[extracted_function_reduction.scala 149:20]
  wire  br_8_io_Out_0_valid; // @[extracted_function_reduction.scala 149:20]
  wire [4:0] br_8_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 149:20]
  wire  br_8_io_Out_0_bits_control; // @[extracted_function_reduction.scala 149:20]
  wire  ret_9_clock; // @[extracted_function_reduction.scala 152:21]
  wire  ret_9_reset; // @[extracted_function_reduction.scala 152:21]
  wire  ret_9_io_In_enable_ready; // @[extracted_function_reduction.scala 152:21]
  wire  ret_9_io_In_enable_valid; // @[extracted_function_reduction.scala 152:21]
  wire [4:0] ret_9_io_In_enable_bits_taskID; // @[extracted_function_reduction.scala 152:21]
  wire  ret_9_io_In_enable_bits_control; // @[extracted_function_reduction.scala 152:21]
  wire  ret_9_io_Out_ready; // @[extracted_function_reduction.scala 152:21]
  wire  ret_9_io_Out_valid; // @[extracted_function_reduction.scala 152:21]
  wire [4:0] ret_9_io_Out_bits_enable_taskID; // @[extracted_function_reduction.scala 152:21]
  wire  ret_9_io_Out_bits_enable_control; // @[extracted_function_reduction.scala 152:21]
  wire  phi_pw_conv_reduction_s1_k_014310_clock; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_reset; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_enable_ready; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_enable_valid; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_enable_bits_control; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_InData_0_ready; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_InData_0_valid; // @[extracted_function_reduction.scala 155:49]
  wire [4:0] phi_pw_conv_reduction_s1_k_014310_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 155:49]
  wire [31:0] phi_pw_conv_reduction_s1_k_014310_io_InData_0_bits_data; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_InData_1_ready; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_InData_1_valid; // @[extracted_function_reduction.scala 155:49]
  wire [4:0] phi_pw_conv_reduction_s1_k_014310_io_InData_1_bits_taskID; // @[extracted_function_reduction.scala 155:49]
  wire [31:0] phi_pw_conv_reduction_s1_k_014310_io_InData_1_bits_data; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_Mask_ready; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_Mask_valid; // @[extracted_function_reduction.scala 155:49]
  wire [1:0] phi_pw_conv_reduction_s1_k_014310_io_Mask_bits; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_Out_0_ready; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_Out_0_valid; // @[extracted_function_reduction.scala 155:49]
  wire [31:0] phi_pw_conv_reduction_s1_k_014310_io_Out_0_bits_data; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_Out_1_ready; // @[extracted_function_reduction.scala 155:49]
  wire  phi_pw_conv_reduction_s1_k_014310_io_Out_1_valid; // @[extracted_function_reduction.scala 155:49]
  wire [31:0] phi_pw_conv_reduction_s1_k_014310_io_Out_1_bits_data; // @[extracted_function_reduction.scala 155:49]
  wire  binaryOp_sub11_clock; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_reset; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_io_enable_ready; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_io_enable_valid; // @[extracted_function_reduction.scala 158:30]
  wire [4:0] binaryOp_sub11_io_enable_bits_taskID; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_io_enable_bits_control; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_io_Out_0_ready; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_io_Out_0_valid; // @[extracted_function_reduction.scala 158:30]
  wire [31:0] binaryOp_sub11_io_Out_0_bits_data; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_io_LeftIO_ready; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_io_LeftIO_valid; // @[extracted_function_reduction.scala 158:30]
  wire [31:0] binaryOp_sub11_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_io_RightIO_ready; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_sub11_io_RightIO_valid; // @[extracted_function_reduction.scala 158:30]
  wire [31:0] binaryOp_sub11_io_RightIO_bits_data; // @[extracted_function_reduction.scala 158:30]
  wire  binaryOp_mul112_clock; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_reset; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_io_enable_ready; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_io_enable_valid; // @[extracted_function_reduction.scala 161:31]
  wire [4:0] binaryOp_mul112_io_enable_bits_taskID; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_io_enable_bits_control; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_io_Out_0_ready; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_io_Out_0_valid; // @[extracted_function_reduction.scala 161:31]
  wire [31:0] binaryOp_mul112_io_Out_0_bits_data; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_io_LeftIO_ready; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_io_LeftIO_valid; // @[extracted_function_reduction.scala 161:31]
  wire [31:0] binaryOp_mul112_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_io_RightIO_ready; // @[extracted_function_reduction.scala 161:31]
  wire  binaryOp_mul112_io_RightIO_valid; // @[extracted_function_reduction.scala 161:31]
  wire [31:0] binaryOp_mul112_io_RightIO_bits_data; // @[extracted_function_reduction.scala 161:31]
  wire  br_13_clock; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_reset; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_enable_ready; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_enable_valid; // @[extracted_function_reduction.scala 164:21]
  wire [4:0] br_13_io_enable_bits_taskID; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_enable_bits_control; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_CmpIO_ready; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_CmpIO_valid; // @[extracted_function_reduction.scala 164:21]
  wire [4:0] br_13_io_CmpIO_bits_taskID; // @[extracted_function_reduction.scala 164:21]
  wire [31:0] br_13_io_CmpIO_bits_data; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_TrueOutput_0_ready; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 164:21]
  wire [4:0] br_13_io_TrueOutput_0_bits_taskID; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_FalseOutput_0_ready; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 164:21]
  wire [4:0] br_13_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 164:21]
  wire  br_13_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 164:21]
  wire  br_14_clock; // @[extracted_function_reduction.scala 167:21]
  wire  br_14_reset; // @[extracted_function_reduction.scala 167:21]
  wire  br_14_io_enable_ready; // @[extracted_function_reduction.scala 167:21]
  wire  br_14_io_enable_valid; // @[extracted_function_reduction.scala 167:21]
  wire [4:0] br_14_io_enable_bits_taskID; // @[extracted_function_reduction.scala 167:21]
  wire  br_14_io_enable_bits_control; // @[extracted_function_reduction.scala 167:21]
  wire  br_14_io_Out_0_ready; // @[extracted_function_reduction.scala 167:21]
  wire  br_14_io_Out_0_valid; // @[extracted_function_reduction.scala 167:21]
  wire [4:0] br_14_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 167:21]
  wire  br_14_io_Out_0_bits_control; // @[extracted_function_reduction.scala 167:21]
  wire  br_15_clock; // @[extracted_function_reduction.scala 170:21]
  wire  br_15_reset; // @[extracted_function_reduction.scala 170:21]
  wire  br_15_io_enable_ready; // @[extracted_function_reduction.scala 170:21]
  wire  br_15_io_enable_valid; // @[extracted_function_reduction.scala 170:21]
  wire [4:0] br_15_io_enable_bits_taskID; // @[extracted_function_reduction.scala 170:21]
  wire  br_15_io_enable_bits_control; // @[extracted_function_reduction.scala 170:21]
  wire  br_15_io_Out_0_ready; // @[extracted_function_reduction.scala 170:21]
  wire  br_15_io_Out_0_valid; // @[extracted_function_reduction.scala 170:21]
  wire [4:0] br_15_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 170:21]
  wire  br_15_io_Out_0_bits_control; // @[extracted_function_reduction.scala 170:21]
  wire  binaryOp_inc6416_clock; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_reset; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_enable_ready; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_enable_valid; // @[extracted_function_reduction.scala 173:32]
  wire [4:0] binaryOp_inc6416_io_enable_bits_taskID; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_enable_bits_control; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_Out_0_ready; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_Out_0_valid; // @[extracted_function_reduction.scala 173:32]
  wire [4:0] binaryOp_inc6416_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 173:32]
  wire [31:0] binaryOp_inc6416_io_Out_0_bits_data; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_Out_1_ready; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_Out_1_valid; // @[extracted_function_reduction.scala 173:32]
  wire [31:0] binaryOp_inc6416_io_Out_1_bits_data; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_LeftIO_ready; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_LeftIO_valid; // @[extracted_function_reduction.scala 173:32]
  wire [31:0] binaryOp_inc6416_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_RightIO_ready; // @[extracted_function_reduction.scala 173:32]
  wire  binaryOp_inc6416_io_RightIO_valid; // @[extracted_function_reduction.scala 173:32]
  wire  icmp_exitcond14817_clock; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_reset; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_io_enable_ready; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_io_enable_valid; // @[extracted_function_reduction.scala 176:34]
  wire [4:0] icmp_exitcond14817_io_enable_bits_taskID; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_io_enable_bits_control; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_io_Out_0_ready; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_io_Out_0_valid; // @[extracted_function_reduction.scala 176:34]
  wire [4:0] icmp_exitcond14817_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 176:34]
  wire [31:0] icmp_exitcond14817_io_Out_0_bits_data; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_io_LeftIO_ready; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_io_LeftIO_valid; // @[extracted_function_reduction.scala 176:34]
  wire [31:0] icmp_exitcond14817_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_io_RightIO_ready; // @[extracted_function_reduction.scala 176:34]
  wire  icmp_exitcond14817_io_RightIO_valid; // @[extracted_function_reduction.scala 176:34]
  wire [31:0] icmp_exitcond14817_io_RightIO_bits_data; // @[extracted_function_reduction.scala 176:34]
  wire  br_18_clock; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_reset; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_enable_ready; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_enable_valid; // @[extracted_function_reduction.scala 179:21]
  wire [4:0] br_18_io_enable_bits_taskID; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_enable_bits_control; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_CmpIO_ready; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_CmpIO_valid; // @[extracted_function_reduction.scala 179:21]
  wire [4:0] br_18_io_CmpIO_bits_taskID; // @[extracted_function_reduction.scala 179:21]
  wire [31:0] br_18_io_CmpIO_bits_data; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_TrueOutput_0_ready; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_FalseOutput_0_ready; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 179:21]
  wire [4:0] br_18_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 179:21]
  wire  br_18_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 179:21]
  wire  phi_pw_conv_reduction_s1_y_014019_clock; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_reset; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_enable_ready; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_enable_valid; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_enable_bits_control; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_InData_0_ready; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_InData_0_valid; // @[extracted_function_reduction.scala 182:49]
  wire [4:0] phi_pw_conv_reduction_s1_y_014019_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 182:49]
  wire [31:0] phi_pw_conv_reduction_s1_y_014019_io_InData_0_bits_data; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_InData_1_ready; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_InData_1_valid; // @[extracted_function_reduction.scala 182:49]
  wire [4:0] phi_pw_conv_reduction_s1_y_014019_io_InData_1_bits_taskID; // @[extracted_function_reduction.scala 182:49]
  wire [31:0] phi_pw_conv_reduction_s1_y_014019_io_InData_1_bits_data; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_Mask_ready; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_Mask_valid; // @[extracted_function_reduction.scala 182:49]
  wire [1:0] phi_pw_conv_reduction_s1_y_014019_io_Mask_bits; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_Out_0_ready; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_Out_0_valid; // @[extracted_function_reduction.scala 182:49]
  wire [31:0] phi_pw_conv_reduction_s1_y_014019_io_Out_0_bits_data; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_Out_1_ready; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_Out_1_valid; // @[extracted_function_reduction.scala 182:49]
  wire [31:0] phi_pw_conv_reduction_s1_y_014019_io_Out_1_bits_data; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_Out_2_ready; // @[extracted_function_reduction.scala 182:49]
  wire  phi_pw_conv_reduction_s1_y_014019_io_Out_2_valid; // @[extracted_function_reduction.scala 182:49]
  wire [31:0] phi_pw_conv_reduction_s1_y_014019_io_Out_2_bits_data; // @[extracted_function_reduction.scala 182:49]
  wire  br_20_clock; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_reset; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_enable_ready; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_enable_valid; // @[extracted_function_reduction.scala 185:21]
  wire [4:0] br_20_io_enable_bits_taskID; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_enable_bits_control; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_CmpIO_ready; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_CmpIO_valid; // @[extracted_function_reduction.scala 185:21]
  wire [4:0] br_20_io_CmpIO_bits_taskID; // @[extracted_function_reduction.scala 185:21]
  wire [31:0] br_20_io_CmpIO_bits_data; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_TrueOutput_0_ready; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 185:21]
  wire [4:0] br_20_io_TrueOutput_0_bits_taskID; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_FalseOutput_0_ready; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 185:21]
  wire [4:0] br_20_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 185:21]
  wire  br_20_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 185:21]
  wire  binaryOp_sub821_clock; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_reset; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_io_enable_ready; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_io_enable_valid; // @[extracted_function_reduction.scala 188:31]
  wire [4:0] binaryOp_sub821_io_enable_bits_taskID; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_io_enable_bits_control; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_io_Out_0_ready; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_io_Out_0_valid; // @[extracted_function_reduction.scala 188:31]
  wire [31:0] binaryOp_sub821_io_Out_0_bits_data; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_io_LeftIO_ready; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_io_LeftIO_valid; // @[extracted_function_reduction.scala 188:31]
  wire [31:0] binaryOp_sub821_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_io_RightIO_ready; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_sub821_io_RightIO_valid; // @[extracted_function_reduction.scala 188:31]
  wire [31:0] binaryOp_sub821_io_RightIO_bits_data; // @[extracted_function_reduction.scala 188:31]
  wire  binaryOp_reass_add22_clock; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_reset; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_io_enable_ready; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_io_enable_valid; // @[extracted_function_reduction.scala 191:36]
  wire [4:0] binaryOp_reass_add22_io_enable_bits_taskID; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_io_enable_bits_control; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_io_Out_0_ready; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_io_Out_0_valid; // @[extracted_function_reduction.scala 191:36]
  wire [31:0] binaryOp_reass_add22_io_Out_0_bits_data; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_io_LeftIO_ready; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_io_LeftIO_valid; // @[extracted_function_reduction.scala 191:36]
  wire [31:0] binaryOp_reass_add22_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_io_RightIO_ready; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_add22_io_RightIO_valid; // @[extracted_function_reduction.scala 191:36]
  wire [31:0] binaryOp_reass_add22_io_RightIO_bits_data; // @[extracted_function_reduction.scala 191:36]
  wire  binaryOp_reass_mul23_clock; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_reset; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_io_enable_ready; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_io_enable_valid; // @[extracted_function_reduction.scala 194:36]
  wire [4:0] binaryOp_reass_mul23_io_enable_bits_taskID; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_io_enable_bits_control; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_io_Out_0_ready; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_io_Out_0_valid; // @[extracted_function_reduction.scala 194:36]
  wire [31:0] binaryOp_reass_mul23_io_Out_0_bits_data; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_io_LeftIO_ready; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_io_LeftIO_valid; // @[extracted_function_reduction.scala 194:36]
  wire [31:0] binaryOp_reass_mul23_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_io_RightIO_ready; // @[extracted_function_reduction.scala 194:36]
  wire  binaryOp_reass_mul23_io_RightIO_valid; // @[extracted_function_reduction.scala 194:36]
  wire [31:0] binaryOp_reass_mul23_io_RightIO_bits_data; // @[extracted_function_reduction.scala 194:36]
  wire  br_24_clock; // @[extracted_function_reduction.scala 197:21]
  wire  br_24_reset; // @[extracted_function_reduction.scala 197:21]
  wire  br_24_io_enable_ready; // @[extracted_function_reduction.scala 197:21]
  wire  br_24_io_enable_valid; // @[extracted_function_reduction.scala 197:21]
  wire [4:0] br_24_io_enable_bits_taskID; // @[extracted_function_reduction.scala 197:21]
  wire  br_24_io_enable_bits_control; // @[extracted_function_reduction.scala 197:21]
  wire  br_24_io_Out_0_ready; // @[extracted_function_reduction.scala 197:21]
  wire  br_24_io_Out_0_valid; // @[extracted_function_reduction.scala 197:21]
  wire [4:0] br_24_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 197:21]
  wire  br_24_io_Out_0_bits_control; // @[extracted_function_reduction.scala 197:21]
  wire  br_25_clock; // @[extracted_function_reduction.scala 200:21]
  wire  br_25_reset; // @[extracted_function_reduction.scala 200:21]
  wire  br_25_io_enable_ready; // @[extracted_function_reduction.scala 200:21]
  wire  br_25_io_enable_valid; // @[extracted_function_reduction.scala 200:21]
  wire [4:0] br_25_io_enable_bits_taskID; // @[extracted_function_reduction.scala 200:21]
  wire  br_25_io_enable_bits_control; // @[extracted_function_reduction.scala 200:21]
  wire  br_25_io_Out_0_ready; // @[extracted_function_reduction.scala 200:21]
  wire  br_25_io_Out_0_valid; // @[extracted_function_reduction.scala 200:21]
  wire [4:0] br_25_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 200:21]
  wire  br_25_io_Out_0_bits_control; // @[extracted_function_reduction.scala 200:21]
  wire  binaryOp_inc6126_clock; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_reset; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_enable_ready; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_enable_valid; // @[extracted_function_reduction.scala 203:32]
  wire [4:0] binaryOp_inc6126_io_enable_bits_taskID; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_enable_bits_control; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_Out_0_ready; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_Out_0_valid; // @[extracted_function_reduction.scala 203:32]
  wire [4:0] binaryOp_inc6126_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 203:32]
  wire [31:0] binaryOp_inc6126_io_Out_0_bits_data; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_Out_1_ready; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_Out_1_valid; // @[extracted_function_reduction.scala 203:32]
  wire [31:0] binaryOp_inc6126_io_Out_1_bits_data; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_LeftIO_ready; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_LeftIO_valid; // @[extracted_function_reduction.scala 203:32]
  wire [31:0] binaryOp_inc6126_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_RightIO_ready; // @[extracted_function_reduction.scala 203:32]
  wire  binaryOp_inc6126_io_RightIO_valid; // @[extracted_function_reduction.scala 203:32]
  wire  icmp_exitcond14727_clock; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_reset; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_io_enable_ready; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_io_enable_valid; // @[extracted_function_reduction.scala 206:34]
  wire [4:0] icmp_exitcond14727_io_enable_bits_taskID; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_io_enable_bits_control; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_io_Out_0_ready; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_io_Out_0_valid; // @[extracted_function_reduction.scala 206:34]
  wire [4:0] icmp_exitcond14727_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 206:34]
  wire [31:0] icmp_exitcond14727_io_Out_0_bits_data; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_io_LeftIO_ready; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_io_LeftIO_valid; // @[extracted_function_reduction.scala 206:34]
  wire [31:0] icmp_exitcond14727_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_io_RightIO_ready; // @[extracted_function_reduction.scala 206:34]
  wire  icmp_exitcond14727_io_RightIO_valid; // @[extracted_function_reduction.scala 206:34]
  wire [31:0] icmp_exitcond14727_io_RightIO_bits_data; // @[extracted_function_reduction.scala 206:34]
  wire  br_28_clock; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_reset; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_enable_ready; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_enable_valid; // @[extracted_function_reduction.scala 209:21]
  wire [4:0] br_28_io_enable_bits_taskID; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_enable_bits_control; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_CmpIO_ready; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_CmpIO_valid; // @[extracted_function_reduction.scala 209:21]
  wire [4:0] br_28_io_CmpIO_bits_taskID; // @[extracted_function_reduction.scala 209:21]
  wire [31:0] br_28_io_CmpIO_bits_data; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_TrueOutput_0_ready; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_FalseOutput_0_ready; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 209:21]
  wire [4:0] br_28_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 209:21]
  wire  br_28_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 209:21]
  wire  phi_pw_conv_reduction_s1_x_013829_clock; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_reset; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_enable_ready; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_enable_valid; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_enable_bits_control; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_InData_0_ready; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_InData_0_valid; // @[extracted_function_reduction.scala 212:49]
  wire [4:0] phi_pw_conv_reduction_s1_x_013829_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 212:49]
  wire [31:0] phi_pw_conv_reduction_s1_x_013829_io_InData_0_bits_data; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_InData_1_ready; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_InData_1_valid; // @[extracted_function_reduction.scala 212:49]
  wire [4:0] phi_pw_conv_reduction_s1_x_013829_io_InData_1_bits_taskID; // @[extracted_function_reduction.scala 212:49]
  wire [31:0] phi_pw_conv_reduction_s1_x_013829_io_InData_1_bits_data; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_Mask_ready; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_Mask_valid; // @[extracted_function_reduction.scala 212:49]
  wire [1:0] phi_pw_conv_reduction_s1_x_013829_io_Mask_bits; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_Out_0_ready; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_Out_0_valid; // @[extracted_function_reduction.scala 212:49]
  wire [31:0] phi_pw_conv_reduction_s1_x_013829_io_Out_0_bits_data; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_Out_1_ready; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_Out_1_valid; // @[extracted_function_reduction.scala 212:49]
  wire [31:0] phi_pw_conv_reduction_s1_x_013829_io_Out_1_bits_data; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_Out_2_ready; // @[extracted_function_reduction.scala 212:49]
  wire  phi_pw_conv_reduction_s1_x_013829_io_Out_2_valid; // @[extracted_function_reduction.scala 212:49]
  wire [31:0] phi_pw_conv_reduction_s1_x_013829_io_Out_2_bits_data; // @[extracted_function_reduction.scala 212:49]
  wire  binaryOp_sub1630_clock; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_reset; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_io_enable_ready; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_io_enable_valid; // @[extracted_function_reduction.scala 215:32]
  wire [4:0] binaryOp_sub1630_io_enable_bits_taskID; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_io_enable_bits_control; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_io_Out_0_ready; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_io_Out_0_valid; // @[extracted_function_reduction.scala 215:32]
  wire [31:0] binaryOp_sub1630_io_Out_0_bits_data; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_io_LeftIO_ready; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_io_LeftIO_valid; // @[extracted_function_reduction.scala 215:32]
  wire [31:0] binaryOp_sub1630_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_io_RightIO_ready; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_sub1630_io_RightIO_valid; // @[extracted_function_reduction.scala 215:32]
  wire [31:0] binaryOp_sub1630_io_RightIO_bits_data; // @[extracted_function_reduction.scala 215:32]
  wire  binaryOp_add1031_clock; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_reset; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_io_enable_ready; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_io_enable_valid; // @[extracted_function_reduction.scala 218:32]
  wire [4:0] binaryOp_add1031_io_enable_bits_taskID; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_io_enable_bits_control; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_io_Out_0_ready; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_io_Out_0_valid; // @[extracted_function_reduction.scala 218:32]
  wire [31:0] binaryOp_add1031_io_Out_0_bits_data; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_io_LeftIO_ready; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_io_LeftIO_valid; // @[extracted_function_reduction.scala 218:32]
  wire [31:0] binaryOp_add1031_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_io_RightIO_ready; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1031_io_RightIO_valid; // @[extracted_function_reduction.scala 218:32]
  wire [31:0] binaryOp_add1031_io_RightIO_bits_data; // @[extracted_function_reduction.scala 218:32]
  wire  binaryOp_add1732_clock; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_reset; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_io_enable_ready; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_io_enable_valid; // @[extracted_function_reduction.scala 221:32]
  wire [4:0] binaryOp_add1732_io_enable_bits_taskID; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_io_enable_bits_control; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_io_Out_0_ready; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_io_Out_0_valid; // @[extracted_function_reduction.scala 221:32]
  wire [31:0] binaryOp_add1732_io_Out_0_bits_data; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_io_LeftIO_ready; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_io_LeftIO_valid; // @[extracted_function_reduction.scala 221:32]
  wire [31:0] binaryOp_add1732_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_io_RightIO_ready; // @[extracted_function_reduction.scala 221:32]
  wire  binaryOp_add1732_io_RightIO_valid; // @[extracted_function_reduction.scala 221:32]
  wire [31:0] binaryOp_add1732_io_RightIO_bits_data; // @[extracted_function_reduction.scala 221:32]
  wire  Gep_arrayidx5033_clock; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_reset; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_enable_ready; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_enable_valid; // @[extracted_function_reduction.scala 224:32]
  wire [4:0] Gep_arrayidx5033_io_enable_bits_taskID; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_enable_bits_control; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_Out_0_ready; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_Out_0_valid; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_Out_0_bits_predicate; // @[extracted_function_reduction.scala 224:32]
  wire [4:0] Gep_arrayidx5033_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 224:32]
  wire [31:0] Gep_arrayidx5033_io_Out_0_bits_data; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_baseAddress_ready; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_baseAddress_valid; // @[extracted_function_reduction.scala 224:32]
  wire [4:0] Gep_arrayidx5033_io_baseAddress_bits_taskID; // @[extracted_function_reduction.scala 224:32]
  wire [31:0] Gep_arrayidx5033_io_baseAddress_bits_data; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_idx_0_ready; // @[extracted_function_reduction.scala 224:32]
  wire  Gep_arrayidx5033_io_idx_0_valid; // @[extracted_function_reduction.scala 224:32]
  wire [31:0] Gep_arrayidx5033_io_idx_0_bits_data; // @[extracted_function_reduction.scala 224:32]
  wire  br_34_clock; // @[extracted_function_reduction.scala 227:21]
  wire  br_34_reset; // @[extracted_function_reduction.scala 227:21]
  wire  br_34_io_enable_ready; // @[extracted_function_reduction.scala 227:21]
  wire  br_34_io_enable_valid; // @[extracted_function_reduction.scala 227:21]
  wire [4:0] br_34_io_enable_bits_taskID; // @[extracted_function_reduction.scala 227:21]
  wire  br_34_io_enable_bits_control; // @[extracted_function_reduction.scala 227:21]
  wire  br_34_io_Out_0_ready; // @[extracted_function_reduction.scala 227:21]
  wire  br_34_io_Out_0_valid; // @[extracted_function_reduction.scala 227:21]
  wire [4:0] br_34_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 227:21]
  wire  br_34_io_Out_0_bits_control; // @[extracted_function_reduction.scala 227:21]
  wire  binaryOp_inc5835_clock; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_reset; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_enable_ready; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_enable_valid; // @[extracted_function_reduction.scala 230:32]
  wire [4:0] binaryOp_inc5835_io_enable_bits_taskID; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_enable_bits_control; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_Out_0_ready; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_Out_0_valid; // @[extracted_function_reduction.scala 230:32]
  wire [4:0] binaryOp_inc5835_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 230:32]
  wire [31:0] binaryOp_inc5835_io_Out_0_bits_data; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_Out_1_ready; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_Out_1_valid; // @[extracted_function_reduction.scala 230:32]
  wire [31:0] binaryOp_inc5835_io_Out_1_bits_data; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_LeftIO_ready; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_LeftIO_valid; // @[extracted_function_reduction.scala 230:32]
  wire [31:0] binaryOp_inc5835_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_RightIO_ready; // @[extracted_function_reduction.scala 230:32]
  wire  binaryOp_inc5835_io_RightIO_valid; // @[extracted_function_reduction.scala 230:32]
  wire  icmp_exitcond14636_clock; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_reset; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_io_enable_ready; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_io_enable_valid; // @[extracted_function_reduction.scala 233:34]
  wire [4:0] icmp_exitcond14636_io_enable_bits_taskID; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_io_enable_bits_control; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_io_Out_0_ready; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_io_Out_0_valid; // @[extracted_function_reduction.scala 233:34]
  wire [4:0] icmp_exitcond14636_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 233:34]
  wire [31:0] icmp_exitcond14636_io_Out_0_bits_data; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_io_LeftIO_ready; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_io_LeftIO_valid; // @[extracted_function_reduction.scala 233:34]
  wire [31:0] icmp_exitcond14636_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_io_RightIO_ready; // @[extracted_function_reduction.scala 233:34]
  wire  icmp_exitcond14636_io_RightIO_valid; // @[extracted_function_reduction.scala 233:34]
  wire [31:0] icmp_exitcond14636_io_RightIO_bits_data; // @[extracted_function_reduction.scala 233:34]
  wire  br_37_clock; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_reset; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_enable_ready; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_enable_valid; // @[extracted_function_reduction.scala 236:21]
  wire [4:0] br_37_io_enable_bits_taskID; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_enable_bits_control; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_CmpIO_ready; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_CmpIO_valid; // @[extracted_function_reduction.scala 236:21]
  wire [4:0] br_37_io_CmpIO_bits_taskID; // @[extracted_function_reduction.scala 236:21]
  wire [31:0] br_37_io_CmpIO_bits_data; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_TrueOutput_0_ready; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_FalseOutput_0_ready; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 236:21]
  wire [4:0] br_37_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 236:21]
  wire  br_37_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 236:21]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_clock; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_reset; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_enable_ready; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_enable_valid; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_enable_bits_control; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_0_ready; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_0_valid; // @[extracted_function_reduction.scala 239:55]
  wire [4:0] phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_ready; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_valid; // @[extracted_function_reduction.scala 239:55]
  wire [4:0] phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_bits_taskID; // @[extracted_function_reduction.scala 239:55]
  wire [31:0] phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_bits_data; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_Mask_ready; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_Mask_valid; // @[extracted_function_reduction.scala 239:55]
  wire [1:0] phi_pw_conv_reduction_s1_r_pw__x_013638_io_Mask_bits; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_0_ready; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_0_valid; // @[extracted_function_reduction.scala 239:55]
  wire [31:0] phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_0_bits_data; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_1_ready; // @[extracted_function_reduction.scala 239:55]
  wire  phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_1_valid; // @[extracted_function_reduction.scala 239:55]
  wire [31:0] phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_1_bits_data; // @[extracted_function_reduction.scala 239:55]
  wire  binaryOp_mul2239_clock; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_reset; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_io_enable_ready; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_io_enable_valid; // @[extracted_function_reduction.scala 242:32]
  wire [4:0] binaryOp_mul2239_io_enable_bits_taskID; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_io_enable_bits_control; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_io_Out_0_ready; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_io_Out_0_valid; // @[extracted_function_reduction.scala 242:32]
  wire [31:0] binaryOp_mul2239_io_Out_0_bits_data; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_io_LeftIO_ready; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_io_LeftIO_valid; // @[extracted_function_reduction.scala 242:32]
  wire [31:0] binaryOp_mul2239_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_io_RightIO_ready; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_mul2239_io_RightIO_valid; // @[extracted_function_reduction.scala 242:32]
  wire [31:0] binaryOp_mul2239_io_RightIO_bits_data; // @[extracted_function_reduction.scala 242:32]
  wire  binaryOp_add2340_clock; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_reset; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_io_enable_ready; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_io_enable_valid; // @[extracted_function_reduction.scala 245:32]
  wire [4:0] binaryOp_add2340_io_enable_bits_taskID; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_io_enable_bits_control; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_io_Out_0_ready; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_io_Out_0_valid; // @[extracted_function_reduction.scala 245:32]
  wire [31:0] binaryOp_add2340_io_Out_0_bits_data; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_io_LeftIO_ready; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_io_LeftIO_valid; // @[extracted_function_reduction.scala 245:32]
  wire [31:0] binaryOp_add2340_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_io_RightIO_ready; // @[extracted_function_reduction.scala 245:32]
  wire  binaryOp_add2340_io_RightIO_valid; // @[extracted_function_reduction.scala 245:32]
  wire [31:0] binaryOp_add2340_io_RightIO_bits_data; // @[extracted_function_reduction.scala 245:32]
  wire  br_41_clock; // @[extracted_function_reduction.scala 248:21]
  wire  br_41_reset; // @[extracted_function_reduction.scala 248:21]
  wire  br_41_io_enable_ready; // @[extracted_function_reduction.scala 248:21]
  wire  br_41_io_enable_valid; // @[extracted_function_reduction.scala 248:21]
  wire [4:0] br_41_io_enable_bits_taskID; // @[extracted_function_reduction.scala 248:21]
  wire  br_41_io_enable_bits_control; // @[extracted_function_reduction.scala 248:21]
  wire  br_41_io_Out_0_ready; // @[extracted_function_reduction.scala 248:21]
  wire  br_41_io_Out_0_valid; // @[extracted_function_reduction.scala 248:21]
  wire [4:0] br_41_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 248:21]
  wire  br_41_io_Out_0_bits_control; // @[extracted_function_reduction.scala 248:21]
  wire  phiadd38_lcssa_lcssa42_clock; // @[extracted_function_reduction.scala 251:38]
  wire  phiadd38_lcssa_lcssa42_reset; // @[extracted_function_reduction.scala 251:38]
  wire  phiadd38_lcssa_lcssa42_io_enable_ready; // @[extracted_function_reduction.scala 251:38]
  wire  phiadd38_lcssa_lcssa42_io_enable_valid; // @[extracted_function_reduction.scala 251:38]
  wire  phiadd38_lcssa_lcssa42_io_enable_bits_control; // @[extracted_function_reduction.scala 251:38]
  wire  phiadd38_lcssa_lcssa42_io_InData_0_ready; // @[extracted_function_reduction.scala 251:38]
  wire  phiadd38_lcssa_lcssa42_io_InData_0_valid; // @[extracted_function_reduction.scala 251:38]
  wire [4:0] phiadd38_lcssa_lcssa42_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 251:38]
  wire [31:0] phiadd38_lcssa_lcssa42_io_InData_0_bits_data; // @[extracted_function_reduction.scala 251:38]
  wire  phiadd38_lcssa_lcssa42_io_Out_0_ready; // @[extracted_function_reduction.scala 251:38]
  wire  phiadd38_lcssa_lcssa42_io_Out_0_valid; // @[extracted_function_reduction.scala 251:38]
  wire [31:0] phiadd38_lcssa_lcssa42_io_Out_0_bits_data; // @[extracted_function_reduction.scala 251:38]
  wire  binaryOp_mul4443_clock; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_reset; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_io_enable_ready; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_io_enable_valid; // @[extracted_function_reduction.scala 254:32]
  wire [4:0] binaryOp_mul4443_io_enable_bits_taskID; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_io_enable_bits_control; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_io_Out_0_ready; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_io_Out_0_valid; // @[extracted_function_reduction.scala 254:32]
  wire [31:0] binaryOp_mul4443_io_Out_0_bits_data; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_io_LeftIO_ready; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_io_LeftIO_valid; // @[extracted_function_reduction.scala 254:32]
  wire [31:0] binaryOp_mul4443_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_io_RightIO_ready; // @[extracted_function_reduction.scala 254:32]
  wire  binaryOp_mul4443_io_RightIO_valid; // @[extracted_function_reduction.scala 254:32]
  wire  sextconv4744_clock; // @[extracted_function_reduction.scala 257:28]
  wire  sextconv4744_reset; // @[extracted_function_reduction.scala 257:28]
  wire  sextconv4744_io_Input_ready; // @[extracted_function_reduction.scala 257:28]
  wire  sextconv4744_io_Input_valid; // @[extracted_function_reduction.scala 257:28]
  wire [31:0] sextconv4744_io_Input_bits_data; // @[extracted_function_reduction.scala 257:28]
  wire  sextconv4744_io_enable_ready; // @[extracted_function_reduction.scala 257:28]
  wire  sextconv4744_io_enable_valid; // @[extracted_function_reduction.scala 257:28]
  wire [4:0] sextconv4744_io_enable_bits_taskID; // @[extracted_function_reduction.scala 257:28]
  wire  sextconv4744_io_Out_0_ready; // @[extracted_function_reduction.scala 257:28]
  wire  sextconv4744_io_Out_0_valid; // @[extracted_function_reduction.scala 257:28]
  wire [31:0] sextconv4744_io_Out_0_bits_data; // @[extracted_function_reduction.scala 257:28]
  wire  ld_45_clock; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_reset; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_enable_ready; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_enable_valid; // @[extracted_function_reduction.scala 260:21]
  wire [4:0] ld_45_io_enable_bits_taskID; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_enable_bits_control; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_Out_0_ready; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_Out_0_valid; // @[extracted_function_reduction.scala 260:21]
  wire [31:0] ld_45_io_Out_0_bits_data; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_GepAddr_ready; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_GepAddr_valid; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_GepAddr_bits_predicate; // @[extracted_function_reduction.scala 260:21]
  wire [4:0] ld_45_io_GepAddr_bits_taskID; // @[extracted_function_reduction.scala 260:21]
  wire [31:0] ld_45_io_GepAddr_bits_data; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_memReq_ready; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_memReq_valid; // @[extracted_function_reduction.scala 260:21]
  wire [31:0] ld_45_io_memReq_bits_address; // @[extracted_function_reduction.scala 260:21]
  wire [4:0] ld_45_io_memReq_bits_taskID; // @[extracted_function_reduction.scala 260:21]
  wire  ld_45_io_memResp_valid; // @[extracted_function_reduction.scala 260:21]
  wire [31:0] ld_45_io_memResp_data; // @[extracted_function_reduction.scala 260:21]
  wire  binaryOp_add5246_clock; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_reset; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_io_enable_ready; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_io_enable_valid; // @[extracted_function_reduction.scala 263:32]
  wire [4:0] binaryOp_add5246_io_enable_bits_taskID; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_io_enable_bits_control; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_io_Out_0_ready; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_io_Out_0_valid; // @[extracted_function_reduction.scala 263:32]
  wire [4:0] binaryOp_add5246_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 263:32]
  wire [31:0] binaryOp_add5246_io_Out_0_bits_data; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_io_LeftIO_ready; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_io_LeftIO_valid; // @[extracted_function_reduction.scala 263:32]
  wire [31:0] binaryOp_add5246_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_io_RightIO_ready; // @[extracted_function_reduction.scala 263:32]
  wire  binaryOp_add5246_io_RightIO_valid; // @[extracted_function_reduction.scala 263:32]
  wire [31:0] binaryOp_add5246_io_RightIO_bits_data; // @[extracted_function_reduction.scala 263:32]
  wire  st_47_clock; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_reset; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_enable_ready; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_enable_valid; // @[extracted_function_reduction.scala 266:21]
  wire [4:0] st_47_io_enable_bits_taskID; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_enable_bits_control; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_GepAddr_ready; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_GepAddr_valid; // @[extracted_function_reduction.scala 266:21]
  wire [4:0] st_47_io_GepAddr_bits_taskID; // @[extracted_function_reduction.scala 266:21]
  wire [31:0] st_47_io_GepAddr_bits_data; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_inData_ready; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_inData_valid; // @[extracted_function_reduction.scala 266:21]
  wire [4:0] st_47_io_inData_bits_taskID; // @[extracted_function_reduction.scala 266:21]
  wire [31:0] st_47_io_inData_bits_data; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_memReq_ready; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_memReq_valid; // @[extracted_function_reduction.scala 266:21]
  wire [21:0] st_47_io_memReq_bits_address; // @[extracted_function_reduction.scala 266:21]
  wire [31:0] st_47_io_memReq_bits_data; // @[extracted_function_reduction.scala 266:21]
  wire [4:0] st_47_io_memReq_bits_taskID; // @[extracted_function_reduction.scala 266:21]
  wire  st_47_io_memResp_valid; // @[extracted_function_reduction.scala 266:21]
  wire  binaryOp_inc5548_clock; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_reset; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_enable_ready; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_enable_valid; // @[extracted_function_reduction.scala 269:32]
  wire [4:0] binaryOp_inc5548_io_enable_bits_taskID; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_enable_bits_control; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_Out_0_ready; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_Out_0_valid; // @[extracted_function_reduction.scala 269:32]
  wire [4:0] binaryOp_inc5548_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 269:32]
  wire [31:0] binaryOp_inc5548_io_Out_0_bits_data; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_Out_1_ready; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_Out_1_valid; // @[extracted_function_reduction.scala 269:32]
  wire [31:0] binaryOp_inc5548_io_Out_1_bits_data; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_LeftIO_ready; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_LeftIO_valid; // @[extracted_function_reduction.scala 269:32]
  wire [31:0] binaryOp_inc5548_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_RightIO_ready; // @[extracted_function_reduction.scala 269:32]
  wire  binaryOp_inc5548_io_RightIO_valid; // @[extracted_function_reduction.scala 269:32]
  wire  icmp_exitcond14549_clock; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_reset; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_io_enable_ready; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_io_enable_valid; // @[extracted_function_reduction.scala 272:34]
  wire [4:0] icmp_exitcond14549_io_enable_bits_taskID; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_io_enable_bits_control; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_io_Out_0_ready; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_io_Out_0_valid; // @[extracted_function_reduction.scala 272:34]
  wire [4:0] icmp_exitcond14549_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 272:34]
  wire [31:0] icmp_exitcond14549_io_Out_0_bits_data; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_io_LeftIO_ready; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_io_LeftIO_valid; // @[extracted_function_reduction.scala 272:34]
  wire [31:0] icmp_exitcond14549_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_io_RightIO_ready; // @[extracted_function_reduction.scala 272:34]
  wire  icmp_exitcond14549_io_RightIO_valid; // @[extracted_function_reduction.scala 272:34]
  wire  br_50_clock; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_reset; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_enable_ready; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_enable_valid; // @[extracted_function_reduction.scala 275:21]
  wire [4:0] br_50_io_enable_bits_taskID; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_enable_bits_control; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_CmpIO_ready; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_CmpIO_valid; // @[extracted_function_reduction.scala 275:21]
  wire [4:0] br_50_io_CmpIO_bits_taskID; // @[extracted_function_reduction.scala 275:21]
  wire [31:0] br_50_io_CmpIO_bits_data; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_TrueOutput_0_ready; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_FalseOutput_0_ready; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 275:21]
  wire [4:0] br_50_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 275:21]
  wire  br_50_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 275:21]
  wire  phi_dw_conv_013551_clock; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_reset; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_enable_ready; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_enable_valid; // @[extracted_function_reduction.scala 278:34]
  wire [4:0] phi_dw_conv_013551_io_enable_bits_taskID; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_enable_bits_control; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_InData_0_ready; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_InData_0_valid; // @[extracted_function_reduction.scala 278:34]
  wire [4:0] phi_dw_conv_013551_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_InData_1_ready; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_InData_1_valid; // @[extracted_function_reduction.scala 278:34]
  wire [4:0] phi_dw_conv_013551_io_InData_1_bits_taskID; // @[extracted_function_reduction.scala 278:34]
  wire [31:0] phi_dw_conv_013551_io_InData_1_bits_data; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_Mask_ready; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_Mask_valid; // @[extracted_function_reduction.scala 278:34]
  wire [1:0] phi_dw_conv_013551_io_Mask_bits; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_Out_0_ready; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_013551_io_Out_0_valid; // @[extracted_function_reduction.scala 278:34]
  wire [4:0] phi_dw_conv_013551_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 278:34]
  wire [31:0] phi_dw_conv_013551_io_Out_0_bits_data; // @[extracted_function_reduction.scala 278:34]
  wire  phi_dw_conv_s1_r_dw__y_013452_clock; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_reset; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_enable_ready; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_enable_valid; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_enable_bits_control; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_InData_0_ready; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_InData_0_valid; // @[extracted_function_reduction.scala 281:45]
  wire [4:0] phi_dw_conv_s1_r_dw__y_013452_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_InData_1_ready; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_InData_1_valid; // @[extracted_function_reduction.scala 281:45]
  wire [4:0] phi_dw_conv_s1_r_dw__y_013452_io_InData_1_bits_taskID; // @[extracted_function_reduction.scala 281:45]
  wire [31:0] phi_dw_conv_s1_r_dw__y_013452_io_InData_1_bits_data; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_Mask_ready; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_Mask_valid; // @[extracted_function_reduction.scala 281:45]
  wire [1:0] phi_dw_conv_s1_r_dw__y_013452_io_Mask_bits; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_Out_0_ready; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_Out_0_valid; // @[extracted_function_reduction.scala 281:45]
  wire [31:0] phi_dw_conv_s1_r_dw__y_013452_io_Out_0_bits_data; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_Out_1_ready; // @[extracted_function_reduction.scala 281:45]
  wire  phi_dw_conv_s1_r_dw__y_013452_io_Out_1_valid; // @[extracted_function_reduction.scala 281:45]
  wire [31:0] phi_dw_conv_s1_r_dw__y_013452_io_Out_1_bits_data; // @[extracted_function_reduction.scala 281:45]
  wire  binaryOp_add2853_clock; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_reset; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_io_enable_ready; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_io_enable_valid; // @[extracted_function_reduction.scala 284:32]
  wire [4:0] binaryOp_add2853_io_enable_bits_taskID; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_io_enable_bits_control; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_io_Out_0_ready; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_io_Out_0_valid; // @[extracted_function_reduction.scala 284:32]
  wire [31:0] binaryOp_add2853_io_Out_0_bits_data; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_io_LeftIO_ready; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_io_LeftIO_valid; // @[extracted_function_reduction.scala 284:32]
  wire [31:0] binaryOp_add2853_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_io_RightIO_ready; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_add2853_io_RightIO_valid; // @[extracted_function_reduction.scala 284:32]
  wire [31:0] binaryOp_add2853_io_RightIO_bits_data; // @[extracted_function_reduction.scala 284:32]
  wire  binaryOp_mul2954_clock; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_reset; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_io_enable_ready; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_io_enable_valid; // @[extracted_function_reduction.scala 287:32]
  wire [4:0] binaryOp_mul2954_io_enable_bits_taskID; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_io_enable_bits_control; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_io_Out_0_ready; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_io_Out_0_valid; // @[extracted_function_reduction.scala 287:32]
  wire [31:0] binaryOp_mul2954_io_Out_0_bits_data; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_io_LeftIO_ready; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_io_LeftIO_valid; // @[extracted_function_reduction.scala 287:32]
  wire [31:0] binaryOp_mul2954_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_io_RightIO_ready; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_mul2954_io_RightIO_valid; // @[extracted_function_reduction.scala 287:32]
  wire [31:0] binaryOp_mul2954_io_RightIO_bits_data; // @[extracted_function_reduction.scala 287:32]
  wire  binaryOp_add3055_clock; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_reset; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_io_enable_ready; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_io_enable_valid; // @[extracted_function_reduction.scala 290:32]
  wire [4:0] binaryOp_add3055_io_enable_bits_taskID; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_io_enable_bits_control; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_io_Out_0_ready; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_io_Out_0_valid; // @[extracted_function_reduction.scala 290:32]
  wire [31:0] binaryOp_add3055_io_Out_0_bits_data; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_io_LeftIO_ready; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_io_LeftIO_valid; // @[extracted_function_reduction.scala 290:32]
  wire [31:0] binaryOp_add3055_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_io_RightIO_ready; // @[extracted_function_reduction.scala 290:32]
  wire  binaryOp_add3055_io_RightIO_valid; // @[extracted_function_reduction.scala 290:32]
  wire [31:0] binaryOp_add3055_io_RightIO_bits_data; // @[extracted_function_reduction.scala 290:32]
  wire  br_56_clock; // @[extracted_function_reduction.scala 293:21]
  wire  br_56_reset; // @[extracted_function_reduction.scala 293:21]
  wire  br_56_io_enable_ready; // @[extracted_function_reduction.scala 293:21]
  wire  br_56_io_enable_valid; // @[extracted_function_reduction.scala 293:21]
  wire [4:0] br_56_io_enable_bits_taskID; // @[extracted_function_reduction.scala 293:21]
  wire  br_56_io_enable_bits_control; // @[extracted_function_reduction.scala 293:21]
  wire  br_56_io_Out_0_ready; // @[extracted_function_reduction.scala 293:21]
  wire  br_56_io_Out_0_valid; // @[extracted_function_reduction.scala 293:21]
  wire [4:0] br_56_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 293:21]
  wire  br_56_io_Out_0_bits_control; // @[extracted_function_reduction.scala 293:21]
  wire  phiadd38_lcssa57_clock; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_reset; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_io_enable_ready; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_io_enable_valid; // @[extracted_function_reduction.scala 296:32]
  wire [4:0] phiadd38_lcssa57_io_enable_bits_taskID; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_io_enable_bits_control; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_io_InData_0_ready; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_io_InData_0_valid; // @[extracted_function_reduction.scala 296:32]
  wire [4:0] phiadd38_lcssa57_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 296:32]
  wire [31:0] phiadd38_lcssa57_io_InData_0_bits_data; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_io_Out_0_ready; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_io_Out_0_valid; // @[extracted_function_reduction.scala 296:32]
  wire [4:0] phiadd38_lcssa57_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 296:32]
  wire [31:0] phiadd38_lcssa57_io_Out_0_bits_data; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_io_Out_1_ready; // @[extracted_function_reduction.scala 296:32]
  wire  phiadd38_lcssa57_io_Out_1_valid; // @[extracted_function_reduction.scala 296:32]
  wire [4:0] phiadd38_lcssa57_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 296:32]
  wire [31:0] phiadd38_lcssa57_io_Out_1_bits_data; // @[extracted_function_reduction.scala 296:32]
  wire  binaryOp_inc4158_clock; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_reset; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_enable_ready; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_enable_valid; // @[extracted_function_reduction.scala 299:32]
  wire [4:0] binaryOp_inc4158_io_enable_bits_taskID; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_enable_bits_control; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_Out_0_ready; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_Out_0_valid; // @[extracted_function_reduction.scala 299:32]
  wire [4:0] binaryOp_inc4158_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 299:32]
  wire [31:0] binaryOp_inc4158_io_Out_0_bits_data; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_Out_1_ready; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_Out_1_valid; // @[extracted_function_reduction.scala 299:32]
  wire [31:0] binaryOp_inc4158_io_Out_1_bits_data; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_LeftIO_ready; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_LeftIO_valid; // @[extracted_function_reduction.scala 299:32]
  wire [31:0] binaryOp_inc4158_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_RightIO_ready; // @[extracted_function_reduction.scala 299:32]
  wire  binaryOp_inc4158_io_RightIO_valid; // @[extracted_function_reduction.scala 299:32]
  wire  icmp_exitcond14459_clock; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_reset; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_io_enable_ready; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_io_enable_valid; // @[extracted_function_reduction.scala 302:34]
  wire [4:0] icmp_exitcond14459_io_enable_bits_taskID; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_io_enable_bits_control; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_io_Out_0_ready; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_io_Out_0_valid; // @[extracted_function_reduction.scala 302:34]
  wire [4:0] icmp_exitcond14459_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 302:34]
  wire [31:0] icmp_exitcond14459_io_Out_0_bits_data; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_io_LeftIO_ready; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_io_LeftIO_valid; // @[extracted_function_reduction.scala 302:34]
  wire [31:0] icmp_exitcond14459_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_io_RightIO_ready; // @[extracted_function_reduction.scala 302:34]
  wire  icmp_exitcond14459_io_RightIO_valid; // @[extracted_function_reduction.scala 302:34]
  wire  br_60_clock; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_reset; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_enable_ready; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_enable_valid; // @[extracted_function_reduction.scala 305:21]
  wire [4:0] br_60_io_enable_bits_taskID; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_enable_bits_control; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_CmpIO_ready; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_CmpIO_valid; // @[extracted_function_reduction.scala 305:21]
  wire [4:0] br_60_io_CmpIO_bits_taskID; // @[extracted_function_reduction.scala 305:21]
  wire [31:0] br_60_io_CmpIO_bits_data; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_TrueOutput_0_ready; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_FalseOutput_0_ready; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 305:21]
  wire [4:0] br_60_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 305:21]
  wire  br_60_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 305:21]
  wire  phi_dw_conv_113361_clock; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_reset; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_enable_ready; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_enable_valid; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_enable_bits_control; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_InData_0_ready; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_InData_0_valid; // @[extracted_function_reduction.scala 308:34]
  wire [4:0] phi_dw_conv_113361_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 308:34]
  wire [31:0] phi_dw_conv_113361_io_InData_0_bits_data; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_InData_1_ready; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_InData_1_valid; // @[extracted_function_reduction.scala 308:34]
  wire [4:0] phi_dw_conv_113361_io_InData_1_bits_taskID; // @[extracted_function_reduction.scala 308:34]
  wire [31:0] phi_dw_conv_113361_io_InData_1_bits_data; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_Mask_ready; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_Mask_valid; // @[extracted_function_reduction.scala 308:34]
  wire [1:0] phi_dw_conv_113361_io_Mask_bits; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_Out_0_ready; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_113361_io_Out_0_valid; // @[extracted_function_reduction.scala 308:34]
  wire [31:0] phi_dw_conv_113361_io_Out_0_bits_data; // @[extracted_function_reduction.scala 308:34]
  wire  phi_dw_conv_s1_r_dw__x_013262_clock; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_reset; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_enable_ready; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_enable_valid; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_enable_bits_control; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_InData_0_ready; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_InData_0_valid; // @[extracted_function_reduction.scala 311:45]
  wire [4:0] phi_dw_conv_s1_r_dw__x_013262_io_InData_0_bits_taskID; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_InData_1_ready; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_InData_1_valid; // @[extracted_function_reduction.scala 311:45]
  wire [4:0] phi_dw_conv_s1_r_dw__x_013262_io_InData_1_bits_taskID; // @[extracted_function_reduction.scala 311:45]
  wire [31:0] phi_dw_conv_s1_r_dw__x_013262_io_InData_1_bits_data; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_Mask_ready; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_Mask_valid; // @[extracted_function_reduction.scala 311:45]
  wire [1:0] phi_dw_conv_s1_r_dw__x_013262_io_Mask_bits; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_Out_0_ready; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_Out_0_valid; // @[extracted_function_reduction.scala 311:45]
  wire [31:0] phi_dw_conv_s1_r_dw__x_013262_io_Out_0_bits_data; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_Out_1_ready; // @[extracted_function_reduction.scala 311:45]
  wire  phi_dw_conv_s1_r_dw__x_013262_io_Out_1_valid; // @[extracted_function_reduction.scala 311:45]
  wire [31:0] phi_dw_conv_s1_r_dw__x_013262_io_Out_1_bits_data; // @[extracted_function_reduction.scala 311:45]
  wire  binaryOp_add3563_clock; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_reset; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_io_enable_ready; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_io_enable_valid; // @[extracted_function_reduction.scala 314:32]
  wire [4:0] binaryOp_add3563_io_enable_bits_taskID; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_io_enable_bits_control; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_io_Out_0_ready; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_io_Out_0_valid; // @[extracted_function_reduction.scala 314:32]
  wire [31:0] binaryOp_add3563_io_Out_0_bits_data; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_io_LeftIO_ready; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_io_LeftIO_valid; // @[extracted_function_reduction.scala 314:32]
  wire [31:0] binaryOp_add3563_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_io_RightIO_ready; // @[extracted_function_reduction.scala 314:32]
  wire  binaryOp_add3563_io_RightIO_valid; // @[extracted_function_reduction.scala 314:32]
  wire [31:0] binaryOp_add3563_io_RightIO_bits_data; // @[extracted_function_reduction.scala 314:32]
  wire  Gep_arrayidx64_clock; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_reset; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_enable_ready; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_enable_valid; // @[extracted_function_reduction.scala 317:30]
  wire [4:0] Gep_arrayidx64_io_enable_bits_taskID; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_enable_bits_control; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_Out_0_ready; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_Out_0_valid; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_Out_0_bits_predicate; // @[extracted_function_reduction.scala 317:30]
  wire [4:0] Gep_arrayidx64_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 317:30]
  wire [31:0] Gep_arrayidx64_io_Out_0_bits_data; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_baseAddress_ready; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_baseAddress_valid; // @[extracted_function_reduction.scala 317:30]
  wire [4:0] Gep_arrayidx64_io_baseAddress_bits_taskID; // @[extracted_function_reduction.scala 317:30]
  wire [31:0] Gep_arrayidx64_io_baseAddress_bits_data; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_idx_0_ready; // @[extracted_function_reduction.scala 317:30]
  wire  Gep_arrayidx64_io_idx_0_valid; // @[extracted_function_reduction.scala 317:30]
  wire [31:0] Gep_arrayidx64_io_idx_0_bits_data; // @[extracted_function_reduction.scala 317:30]
  wire  ld_65_clock; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_reset; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_enable_ready; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_enable_valid; // @[extracted_function_reduction.scala 320:21]
  wire [4:0] ld_65_io_enable_bits_taskID; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_enable_bits_control; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_Out_0_ready; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_Out_0_valid; // @[extracted_function_reduction.scala 320:21]
  wire [31:0] ld_65_io_Out_0_bits_data; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_GepAddr_ready; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_GepAddr_valid; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_GepAddr_bits_predicate; // @[extracted_function_reduction.scala 320:21]
  wire [4:0] ld_65_io_GepAddr_bits_taskID; // @[extracted_function_reduction.scala 320:21]
  wire [31:0] ld_65_io_GepAddr_bits_data; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_memReq_ready; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_memReq_valid; // @[extracted_function_reduction.scala 320:21]
  wire [31:0] ld_65_io_memReq_bits_address; // @[extracted_function_reduction.scala 320:21]
  wire [4:0] ld_65_io_memReq_bits_taskID; // @[extracted_function_reduction.scala 320:21]
  wire  ld_65_io_memResp_valid; // @[extracted_function_reduction.scala 320:21]
  wire [31:0] ld_65_io_memResp_data; // @[extracted_function_reduction.scala 320:21]
  wire  sextconv3766_clock; // @[extracted_function_reduction.scala 323:28]
  wire  sextconv3766_reset; // @[extracted_function_reduction.scala 323:28]
  wire  sextconv3766_io_Input_ready; // @[extracted_function_reduction.scala 323:28]
  wire  sextconv3766_io_Input_valid; // @[extracted_function_reduction.scala 323:28]
  wire [31:0] sextconv3766_io_Input_bits_data; // @[extracted_function_reduction.scala 323:28]
  wire  sextconv3766_io_enable_ready; // @[extracted_function_reduction.scala 323:28]
  wire  sextconv3766_io_enable_valid; // @[extracted_function_reduction.scala 323:28]
  wire [4:0] sextconv3766_io_enable_bits_taskID; // @[extracted_function_reduction.scala 323:28]
  wire  sextconv3766_io_Out_0_ready; // @[extracted_function_reduction.scala 323:28]
  wire  sextconv3766_io_Out_0_valid; // @[extracted_function_reduction.scala 323:28]
  wire [31:0] sextconv3766_io_Out_0_bits_data; // @[extracted_function_reduction.scala 323:28]
  wire  binaryOp_add3867_clock; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_reset; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_enable_ready; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_enable_valid; // @[extracted_function_reduction.scala 326:32]
  wire [4:0] binaryOp_add3867_io_enable_bits_taskID; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_enable_bits_control; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_Out_0_ready; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_Out_0_valid; // @[extracted_function_reduction.scala 326:32]
  wire [4:0] binaryOp_add3867_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 326:32]
  wire [31:0] binaryOp_add3867_io_Out_0_bits_data; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_Out_1_ready; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_Out_1_valid; // @[extracted_function_reduction.scala 326:32]
  wire [4:0] binaryOp_add3867_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 326:32]
  wire [31:0] binaryOp_add3867_io_Out_1_bits_data; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_LeftIO_ready; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_LeftIO_valid; // @[extracted_function_reduction.scala 326:32]
  wire [31:0] binaryOp_add3867_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_RightIO_ready; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_add3867_io_RightIO_valid; // @[extracted_function_reduction.scala 326:32]
  wire [31:0] binaryOp_add3867_io_RightIO_bits_data; // @[extracted_function_reduction.scala 326:32]
  wire  binaryOp_inc68_clock; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_reset; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_enable_ready; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_enable_valid; // @[extracted_function_reduction.scala 329:30]
  wire [4:0] binaryOp_inc68_io_enable_bits_taskID; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_enable_bits_control; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_Out_0_ready; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_Out_0_valid; // @[extracted_function_reduction.scala 329:30]
  wire [4:0] binaryOp_inc68_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 329:30]
  wire [31:0] binaryOp_inc68_io_Out_0_bits_data; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_Out_1_ready; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_Out_1_valid; // @[extracted_function_reduction.scala 329:30]
  wire [31:0] binaryOp_inc68_io_Out_1_bits_data; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_LeftIO_ready; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_LeftIO_valid; // @[extracted_function_reduction.scala 329:30]
  wire [31:0] binaryOp_inc68_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_RightIO_ready; // @[extracted_function_reduction.scala 329:30]
  wire  binaryOp_inc68_io_RightIO_valid; // @[extracted_function_reduction.scala 329:30]
  wire  icmp_exitcond69_clock; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_reset; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_io_enable_ready; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_io_enable_valid; // @[extracted_function_reduction.scala 332:31]
  wire [4:0] icmp_exitcond69_io_enable_bits_taskID; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_io_enable_bits_control; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_io_Out_0_ready; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_io_Out_0_valid; // @[extracted_function_reduction.scala 332:31]
  wire [4:0] icmp_exitcond69_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 332:31]
  wire [31:0] icmp_exitcond69_io_Out_0_bits_data; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_io_LeftIO_ready; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_io_LeftIO_valid; // @[extracted_function_reduction.scala 332:31]
  wire [31:0] icmp_exitcond69_io_LeftIO_bits_data; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_io_RightIO_ready; // @[extracted_function_reduction.scala 332:31]
  wire  icmp_exitcond69_io_RightIO_valid; // @[extracted_function_reduction.scala 332:31]
  wire  br_70_clock; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_reset; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_enable_ready; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_enable_valid; // @[extracted_function_reduction.scala 335:21]
  wire [4:0] br_70_io_enable_bits_taskID; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_enable_bits_control; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_CmpIO_ready; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_CmpIO_valid; // @[extracted_function_reduction.scala 335:21]
  wire [4:0] br_70_io_CmpIO_bits_taskID; // @[extracted_function_reduction.scala 335:21]
  wire [31:0] br_70_io_CmpIO_bits_data; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_TrueOutput_0_ready; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_FalseOutput_0_ready; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 335:21]
  wire [4:0] br_70_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 335:21]
  wire  br_70_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 335:21]
  wire  const0_clock; // @[extracted_function_reduction.scala 344:22]
  wire  const0_reset; // @[extracted_function_reduction.scala 344:22]
  wire  const0_io_enable_ready; // @[extracted_function_reduction.scala 344:22]
  wire  const0_io_enable_valid; // @[extracted_function_reduction.scala 344:22]
  wire [4:0] const0_io_enable_bits_taskID; // @[extracted_function_reduction.scala 344:22]
  wire  const0_io_Out_ready; // @[extracted_function_reduction.scala 344:22]
  wire  const0_io_Out_valid; // @[extracted_function_reduction.scala 344:22]
  wire  const1_clock; // @[extracted_function_reduction.scala 347:22]
  wire  const1_reset; // @[extracted_function_reduction.scala 347:22]
  wire  const1_io_enable_ready; // @[extracted_function_reduction.scala 347:22]
  wire  const1_io_enable_valid; // @[extracted_function_reduction.scala 347:22]
  wire [4:0] const1_io_enable_bits_taskID; // @[extracted_function_reduction.scala 347:22]
  wire  const1_io_Out_ready; // @[extracted_function_reduction.scala 347:22]
  wire  const1_io_Out_valid; // @[extracted_function_reduction.scala 347:22]
  wire  const2_clock; // @[extracted_function_reduction.scala 350:22]
  wire  const2_reset; // @[extracted_function_reduction.scala 350:22]
  wire  const2_io_enable_ready; // @[extracted_function_reduction.scala 350:22]
  wire  const2_io_enable_valid; // @[extracted_function_reduction.scala 350:22]
  wire [4:0] const2_io_enable_bits_taskID; // @[extracted_function_reduction.scala 350:22]
  wire  const2_io_Out_ready; // @[extracted_function_reduction.scala 350:22]
  wire  const2_io_Out_valid; // @[extracted_function_reduction.scala 350:22]
  wire  const3_clock; // @[extracted_function_reduction.scala 353:22]
  wire  const3_reset; // @[extracted_function_reduction.scala 353:22]
  wire  const3_io_enable_ready; // @[extracted_function_reduction.scala 353:22]
  wire  const3_io_enable_valid; // @[extracted_function_reduction.scala 353:22]
  wire [4:0] const3_io_enable_bits_taskID; // @[extracted_function_reduction.scala 353:22]
  wire  const3_io_Out_ready; // @[extracted_function_reduction.scala 353:22]
  wire  const3_io_Out_valid; // @[extracted_function_reduction.scala 353:22]
  wire [4:0] const3_io_Out_bits_taskID; // @[extracted_function_reduction.scala 353:22]
  wire  const4_clock; // @[extracted_function_reduction.scala 356:22]
  wire  const4_reset; // @[extracted_function_reduction.scala 356:22]
  wire  const4_io_enable_ready; // @[extracted_function_reduction.scala 356:22]
  wire  const4_io_enable_valid; // @[extracted_function_reduction.scala 356:22]
  wire [4:0] const4_io_enable_bits_taskID; // @[extracted_function_reduction.scala 356:22]
  wire  const4_io_Out_ready; // @[extracted_function_reduction.scala 356:22]
  wire  const4_io_Out_valid; // @[extracted_function_reduction.scala 356:22]
  wire  const5_clock; // @[extracted_function_reduction.scala 359:22]
  wire  const5_reset; // @[extracted_function_reduction.scala 359:22]
  wire  const5_io_enable_ready; // @[extracted_function_reduction.scala 359:22]
  wire  const5_io_enable_valid; // @[extracted_function_reduction.scala 359:22]
  wire [4:0] const5_io_enable_bits_taskID; // @[extracted_function_reduction.scala 359:22]
  wire  const5_io_Out_ready; // @[extracted_function_reduction.scala 359:22]
  wire  const5_io_Out_valid; // @[extracted_function_reduction.scala 359:22]
  wire  const6_clock; // @[extracted_function_reduction.scala 362:22]
  wire  const6_reset; // @[extracted_function_reduction.scala 362:22]
  wire  const6_io_enable_ready; // @[extracted_function_reduction.scala 362:22]
  wire  const6_io_enable_valid; // @[extracted_function_reduction.scala 362:22]
  wire [4:0] const6_io_enable_bits_taskID; // @[extracted_function_reduction.scala 362:22]
  wire  const6_io_Out_ready; // @[extracted_function_reduction.scala 362:22]
  wire  const6_io_Out_valid; // @[extracted_function_reduction.scala 362:22]
  wire  const7_clock; // @[extracted_function_reduction.scala 365:22]
  wire  const7_reset; // @[extracted_function_reduction.scala 365:22]
  wire  const7_io_enable_ready; // @[extracted_function_reduction.scala 365:22]
  wire  const7_io_enable_valid; // @[extracted_function_reduction.scala 365:22]
  wire [4:0] const7_io_enable_bits_taskID; // @[extracted_function_reduction.scala 365:22]
  wire  const7_io_Out_ready; // @[extracted_function_reduction.scala 365:22]
  wire  const7_io_Out_valid; // @[extracted_function_reduction.scala 365:22]
  wire [4:0] const7_io_Out_bits_taskID; // @[extracted_function_reduction.scala 365:22]
  wire  const8_clock; // @[extracted_function_reduction.scala 368:22]
  wire  const8_reset; // @[extracted_function_reduction.scala 368:22]
  wire  const8_io_enable_ready; // @[extracted_function_reduction.scala 368:22]
  wire  const8_io_enable_valid; // @[extracted_function_reduction.scala 368:22]
  wire [4:0] const8_io_enable_bits_taskID; // @[extracted_function_reduction.scala 368:22]
  wire  const8_io_Out_ready; // @[extracted_function_reduction.scala 368:22]
  wire  const8_io_Out_valid; // @[extracted_function_reduction.scala 368:22]
  wire [4:0] const8_io_Out_bits_taskID; // @[extracted_function_reduction.scala 368:22]
  wire  const9_clock; // @[extracted_function_reduction.scala 371:22]
  wire  const9_reset; // @[extracted_function_reduction.scala 371:22]
  wire  const9_io_enable_ready; // @[extracted_function_reduction.scala 371:22]
  wire  const9_io_enable_valid; // @[extracted_function_reduction.scala 371:22]
  wire [4:0] const9_io_enable_bits_taskID; // @[extracted_function_reduction.scala 371:22]
  wire  const9_io_Out_ready; // @[extracted_function_reduction.scala 371:22]
  wire  const9_io_Out_valid; // @[extracted_function_reduction.scala 371:22]
  wire  const10_clock; // @[extracted_function_reduction.scala 374:23]
  wire  const10_reset; // @[extracted_function_reduction.scala 374:23]
  wire  const10_io_enable_ready; // @[extracted_function_reduction.scala 374:23]
  wire  const10_io_enable_valid; // @[extracted_function_reduction.scala 374:23]
  wire [4:0] const10_io_enable_bits_taskID; // @[extracted_function_reduction.scala 374:23]
  wire  const10_io_Out_ready; // @[extracted_function_reduction.scala 374:23]
  wire  const10_io_Out_valid; // @[extracted_function_reduction.scala 374:23]
  wire  const11_clock; // @[extracted_function_reduction.scala 377:23]
  wire  const11_reset; // @[extracted_function_reduction.scala 377:23]
  wire  const11_io_enable_ready; // @[extracted_function_reduction.scala 377:23]
  wire  const11_io_enable_valid; // @[extracted_function_reduction.scala 377:23]
  wire [4:0] const11_io_enable_bits_taskID; // @[extracted_function_reduction.scala 377:23]
  wire  const11_io_Out_ready; // @[extracted_function_reduction.scala 377:23]
  wire  const11_io_Out_valid; // @[extracted_function_reduction.scala 377:23]
  wire [4:0] const11_io_Out_bits_taskID; // @[extracted_function_reduction.scala 377:23]
  wire  const12_clock; // @[extracted_function_reduction.scala 380:23]
  wire  const12_reset; // @[extracted_function_reduction.scala 380:23]
  wire  const12_io_enable_ready; // @[extracted_function_reduction.scala 380:23]
  wire  const12_io_enable_valid; // @[extracted_function_reduction.scala 380:23]
  wire [4:0] const12_io_enable_bits_taskID; // @[extracted_function_reduction.scala 380:23]
  wire  const12_io_Out_ready; // @[extracted_function_reduction.scala 380:23]
  wire  const12_io_Out_valid; // @[extracted_function_reduction.scala 380:23]
  wire  const13_clock; // @[extracted_function_reduction.scala 383:23]
  wire  const13_reset; // @[extracted_function_reduction.scala 383:23]
  wire  const13_io_enable_ready; // @[extracted_function_reduction.scala 383:23]
  wire  const13_io_enable_valid; // @[extracted_function_reduction.scala 383:23]
  wire [4:0] const13_io_enable_bits_taskID; // @[extracted_function_reduction.scala 383:23]
  wire  const13_io_Out_ready; // @[extracted_function_reduction.scala 383:23]
  wire  const13_io_Out_valid; // @[extracted_function_reduction.scala 383:23]
  UnifiedController MemCtrl ( // @[extracted_function_reduction.scala 45:23]
    .clock(MemCtrl_clock),
    .reset(MemCtrl_reset),
    .io_WriteIn_0_ready(MemCtrl_io_WriteIn_0_ready),
    .io_WriteIn_0_valid(MemCtrl_io_WriteIn_0_valid),
    .io_WriteIn_0_bits_address(MemCtrl_io_WriteIn_0_bits_address),
    .io_WriteIn_0_bits_data(MemCtrl_io_WriteIn_0_bits_data),
    .io_WriteIn_0_bits_taskID(MemCtrl_io_WriteIn_0_bits_taskID),
    .io_WriteOut_0_valid(MemCtrl_io_WriteOut_0_valid),
    .io_ReadIn_0_ready(MemCtrl_io_ReadIn_0_ready),
    .io_ReadIn_0_valid(MemCtrl_io_ReadIn_0_valid),
    .io_ReadIn_0_bits_address(MemCtrl_io_ReadIn_0_bits_address),
    .io_ReadIn_0_bits_taskID(MemCtrl_io_ReadIn_0_bits_taskID),
    .io_ReadIn_1_ready(MemCtrl_io_ReadIn_1_ready),
    .io_ReadIn_1_valid(MemCtrl_io_ReadIn_1_valid),
    .io_ReadIn_1_bits_address(MemCtrl_io_ReadIn_1_bits_address),
    .io_ReadIn_1_bits_taskID(MemCtrl_io_ReadIn_1_bits_taskID),
    .io_ReadOut_0_valid(MemCtrl_io_ReadOut_0_valid),
    .io_ReadOut_0_data(MemCtrl_io_ReadOut_0_data),
    .io_ReadOut_1_valid(MemCtrl_io_ReadOut_1_valid),
    .io_ReadOut_1_data(MemCtrl_io_ReadOut_1_data),
    .io_MemResp_valid(MemCtrl_io_MemResp_valid),
    .io_MemResp_bits_data(MemCtrl_io_MemResp_bits_data),
    .io_MemResp_bits_tag(MemCtrl_io_MemResp_bits_tag),
    .io_MemResp_bits_iswrite(MemCtrl_io_MemResp_bits_iswrite),
    .io_MemReq_ready(MemCtrl_io_MemReq_ready),
    .io_MemReq_valid(MemCtrl_io_MemReq_valid),
    .io_MemReq_bits_addr(MemCtrl_io_MemReq_bits_addr),
    .io_MemReq_bits_data(MemCtrl_io_MemReq_bits_data),
    .io_MemReq_bits_mask(MemCtrl_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(MemCtrl_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(MemCtrl_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(MemCtrl_io_MemReq_bits_iswrite)
  );
  SplitCallNew InputSplitter ( // @[extracted_function_reduction.scala 53:29]
    .clock(InputSplitter_clock),
    .reset(InputSplitter_reset),
    .io_In_ready(InputSplitter_io_In_ready),
    .io_In_valid(InputSplitter_io_In_valid),
    .io_In_bits_enable_taskID(InputSplitter_io_In_bits_enable_taskID),
    .io_In_bits_enable_control(InputSplitter_io_In_bits_enable_control),
    .io_In_bits_data_field10_data(InputSplitter_io_In_bits_data_field10_data),
    .io_In_bits_data_field9_data(InputSplitter_io_In_bits_data_field9_data),
    .io_In_bits_data_field8_taskID(InputSplitter_io_In_bits_data_field8_taskID),
    .io_In_bits_data_field8_data(InputSplitter_io_In_bits_data_field8_data),
    .io_In_bits_data_field7_data(InputSplitter_io_In_bits_data_field7_data),
    .io_In_bits_data_field6_taskID(InputSplitter_io_In_bits_data_field6_taskID),
    .io_In_bits_data_field6_data(InputSplitter_io_In_bits_data_field6_data),
    .io_In_bits_data_field5_data(InputSplitter_io_In_bits_data_field5_data),
    .io_In_bits_data_field4_taskID(InputSplitter_io_In_bits_data_field4_taskID),
    .io_In_bits_data_field4_data(InputSplitter_io_In_bits_data_field4_data),
    .io_In_bits_data_field3_data(InputSplitter_io_In_bits_data_field3_data),
    .io_In_bits_data_field2_data(InputSplitter_io_In_bits_data_field2_data),
    .io_In_bits_data_field1_taskID(InputSplitter_io_In_bits_data_field1_taskID),
    .io_In_bits_data_field1_data(InputSplitter_io_In_bits_data_field1_data),
    .io_In_bits_data_field0_taskID(InputSplitter_io_In_bits_data_field0_taskID),
    .io_In_bits_data_field0_data(InputSplitter_io_In_bits_data_field0_data),
    .io_Out_enable_ready(InputSplitter_io_Out_enable_ready),
    .io_Out_enable_valid(InputSplitter_io_Out_enable_valid),
    .io_Out_enable_bits_taskID(InputSplitter_io_Out_enable_bits_taskID),
    .io_Out_enable_bits_control(InputSplitter_io_Out_enable_bits_control),
    .io_Out_data_field10_0_ready(InputSplitter_io_Out_data_field10_0_ready),
    .io_Out_data_field10_0_valid(InputSplitter_io_Out_data_field10_0_valid),
    .io_Out_data_field10_0_bits_data(InputSplitter_io_Out_data_field10_0_bits_data),
    .io_Out_data_field9_0_ready(InputSplitter_io_Out_data_field9_0_ready),
    .io_Out_data_field9_0_valid(InputSplitter_io_Out_data_field9_0_valid),
    .io_Out_data_field9_0_bits_data(InputSplitter_io_Out_data_field9_0_bits_data),
    .io_Out_data_field8_0_ready(InputSplitter_io_Out_data_field8_0_ready),
    .io_Out_data_field8_0_valid(InputSplitter_io_Out_data_field8_0_valid),
    .io_Out_data_field8_0_bits_taskID(InputSplitter_io_Out_data_field8_0_bits_taskID),
    .io_Out_data_field8_0_bits_data(InputSplitter_io_Out_data_field8_0_bits_data),
    .io_Out_data_field8_1_ready(InputSplitter_io_Out_data_field8_1_ready),
    .io_Out_data_field8_1_valid(InputSplitter_io_Out_data_field8_1_valid),
    .io_Out_data_field8_1_bits_data(InputSplitter_io_Out_data_field8_1_bits_data),
    .io_Out_data_field8_2_ready(InputSplitter_io_Out_data_field8_2_ready),
    .io_Out_data_field8_2_valid(InputSplitter_io_Out_data_field8_2_valid),
    .io_Out_data_field8_2_bits_data(InputSplitter_io_Out_data_field8_2_bits_data),
    .io_Out_data_field7_0_ready(InputSplitter_io_Out_data_field7_0_ready),
    .io_Out_data_field7_0_valid(InputSplitter_io_Out_data_field7_0_valid),
    .io_Out_data_field7_0_bits_data(InputSplitter_io_Out_data_field7_0_bits_data),
    .io_Out_data_field7_1_ready(InputSplitter_io_Out_data_field7_1_ready),
    .io_Out_data_field7_1_valid(InputSplitter_io_Out_data_field7_1_valid),
    .io_Out_data_field7_1_bits_data(InputSplitter_io_Out_data_field7_1_bits_data),
    .io_Out_data_field6_0_ready(InputSplitter_io_Out_data_field6_0_ready),
    .io_Out_data_field6_0_valid(InputSplitter_io_Out_data_field6_0_valid),
    .io_Out_data_field6_0_bits_taskID(InputSplitter_io_Out_data_field6_0_bits_taskID),
    .io_Out_data_field6_0_bits_data(InputSplitter_io_Out_data_field6_0_bits_data),
    .io_Out_data_field6_1_ready(InputSplitter_io_Out_data_field6_1_ready),
    .io_Out_data_field6_1_valid(InputSplitter_io_Out_data_field6_1_valid),
    .io_Out_data_field6_1_bits_data(InputSplitter_io_Out_data_field6_1_bits_data),
    .io_Out_data_field6_2_ready(InputSplitter_io_Out_data_field6_2_ready),
    .io_Out_data_field6_2_valid(InputSplitter_io_Out_data_field6_2_valid),
    .io_Out_data_field6_2_bits_data(InputSplitter_io_Out_data_field6_2_bits_data),
    .io_Out_data_field5_0_ready(InputSplitter_io_Out_data_field5_0_ready),
    .io_Out_data_field5_0_valid(InputSplitter_io_Out_data_field5_0_valid),
    .io_Out_data_field5_0_bits_data(InputSplitter_io_Out_data_field5_0_bits_data),
    .io_Out_data_field5_1_ready(InputSplitter_io_Out_data_field5_1_ready),
    .io_Out_data_field5_1_valid(InputSplitter_io_Out_data_field5_1_valid),
    .io_Out_data_field5_1_bits_data(InputSplitter_io_Out_data_field5_1_bits_data),
    .io_Out_data_field4_0_ready(InputSplitter_io_Out_data_field4_0_ready),
    .io_Out_data_field4_0_valid(InputSplitter_io_Out_data_field4_0_valid),
    .io_Out_data_field4_0_bits_taskID(InputSplitter_io_Out_data_field4_0_bits_taskID),
    .io_Out_data_field4_0_bits_data(InputSplitter_io_Out_data_field4_0_bits_data),
    .io_Out_data_field4_1_ready(InputSplitter_io_Out_data_field4_1_ready),
    .io_Out_data_field4_1_valid(InputSplitter_io_Out_data_field4_1_valid),
    .io_Out_data_field4_1_bits_data(InputSplitter_io_Out_data_field4_1_bits_data),
    .io_Out_data_field4_2_ready(InputSplitter_io_Out_data_field4_2_ready),
    .io_Out_data_field4_2_valid(InputSplitter_io_Out_data_field4_2_valid),
    .io_Out_data_field4_2_bits_data(InputSplitter_io_Out_data_field4_2_bits_data),
    .io_Out_data_field3_0_ready(InputSplitter_io_Out_data_field3_0_ready),
    .io_Out_data_field3_0_valid(InputSplitter_io_Out_data_field3_0_valid),
    .io_Out_data_field3_0_bits_data(InputSplitter_io_Out_data_field3_0_bits_data),
    .io_Out_data_field2_0_ready(InputSplitter_io_Out_data_field2_0_ready),
    .io_Out_data_field2_0_valid(InputSplitter_io_Out_data_field2_0_valid),
    .io_Out_data_field2_0_bits_data(InputSplitter_io_Out_data_field2_0_bits_data),
    .io_Out_data_field1_0_ready(InputSplitter_io_Out_data_field1_0_ready),
    .io_Out_data_field1_0_valid(InputSplitter_io_Out_data_field1_0_valid),
    .io_Out_data_field1_0_bits_taskID(InputSplitter_io_Out_data_field1_0_bits_taskID),
    .io_Out_data_field1_0_bits_data(InputSplitter_io_Out_data_field1_0_bits_data),
    .io_Out_data_field0_0_ready(InputSplitter_io_Out_data_field0_0_ready),
    .io_Out_data_field0_0_valid(InputSplitter_io_Out_data_field0_0_valid),
    .io_Out_data_field0_0_bits_taskID(InputSplitter_io_Out_data_field0_0_bits_taskID),
    .io_Out_data_field0_0_bits_data(InputSplitter_io_Out_data_field0_0_bits_data)
  );
  LoopBlockNode Loop_0 ( // @[extracted_function_reduction.scala 62:22]
    .clock(Loop_0_clock),
    .reset(Loop_0_reset),
    .io_enable_ready(Loop_0_io_enable_ready),
    .io_enable_valid(Loop_0_io_enable_valid),
    .io_enable_bits_taskID(Loop_0_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_0_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_0_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_0_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_taskID(Loop_0_io_InLiveIn_0_bits_taskID),
    .io_InLiveIn_0_bits_data(Loop_0_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_0_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_0_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_0_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_0_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_0_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_taskID(Loop_0_io_InLiveIn_2_bits_taskID),
    .io_InLiveIn_2_bits_data(Loop_0_io_InLiveIn_2_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_0_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_0_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_taskID(Loop_0_io_OutLiveIn_field2_0_bits_taskID),
    .io_OutLiveIn_field2_0_bits_data(Loop_0_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_0_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_0_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_0_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_0_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_0_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_taskID(Loop_0_io_OutLiveIn_field0_0_bits_taskID),
    .io_OutLiveIn_field0_0_bits_data(Loop_0_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_0_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_0_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_0_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_0_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_0_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_0_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_0_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_0_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_0_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_0_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_0_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_0_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_0_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_0_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_0_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_0_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_0_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_0_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_0_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenIn_1_ready(Loop_0_io_CarryDepenIn_1_ready),
    .io_CarryDepenIn_1_valid(Loop_0_io_CarryDepenIn_1_valid),
    .io_CarryDepenIn_1_bits_taskID(Loop_0_io_CarryDepenIn_1_bits_taskID),
    .io_CarryDepenIn_1_bits_data(Loop_0_io_CarryDepenIn_1_bits_data),
    .io_CarryDepenOut_field1_0_ready(Loop_0_io_CarryDepenOut_field1_0_ready),
    .io_CarryDepenOut_field1_0_valid(Loop_0_io_CarryDepenOut_field1_0_valid),
    .io_CarryDepenOut_field1_0_bits_taskID(Loop_0_io_CarryDepenOut_field1_0_bits_taskID),
    .io_CarryDepenOut_field1_0_bits_data(Loop_0_io_CarryDepenOut_field1_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_0_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_0_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_0_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_0_io_CarryDepenOut_field0_0_bits_data),
    .io_InLiveOut_0_ready(Loop_0_io_InLiveOut_0_ready),
    .io_InLiveOut_0_valid(Loop_0_io_InLiveOut_0_valid),
    .io_InLiveOut_0_bits_taskID(Loop_0_io_InLiveOut_0_bits_taskID),
    .io_InLiveOut_0_bits_data(Loop_0_io_InLiveOut_0_bits_data),
    .io_OutLiveOut_field0_0_ready(Loop_0_io_OutLiveOut_field0_0_ready),
    .io_OutLiveOut_field0_0_valid(Loop_0_io_OutLiveOut_field0_0_valid),
    .io_OutLiveOut_field0_0_bits_taskID(Loop_0_io_OutLiveOut_field0_0_bits_taskID),
    .io_OutLiveOut_field0_0_bits_data(Loop_0_io_OutLiveOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_0_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_0_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_0_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_0_io_loopExit_0_bits_control)
  );
  LoopBlockNode_1 Loop_1 ( // @[extracted_function_reduction.scala 64:22]
    .clock(Loop_1_clock),
    .reset(Loop_1_reset),
    .io_enable_ready(Loop_1_io_enable_ready),
    .io_enable_valid(Loop_1_io_enable_valid),
    .io_enable_bits_taskID(Loop_1_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_1_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_1_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_1_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_1_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_1_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_1_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_taskID(Loop_1_io_InLiveIn_1_bits_taskID),
    .io_InLiveIn_1_bits_data(Loop_1_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_1_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_1_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_1_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_1_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_1_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_data(Loop_1_io_InLiveIn_3_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_1_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_1_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_data(Loop_1_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_1_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_1_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_1_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_1_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_1_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_taskID(Loop_1_io_OutLiveIn_field1_0_bits_taskID),
    .io_OutLiveIn_field1_0_bits_data(Loop_1_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_1_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_1_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_1_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_1_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_1_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_1_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_1_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_1_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_1_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_1_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_1_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_1_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_1_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_1_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_1_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_1_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_1_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_1_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_1_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_1_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_1_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_1_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenIn_1_ready(Loop_1_io_CarryDepenIn_1_ready),
    .io_CarryDepenIn_1_valid(Loop_1_io_CarryDepenIn_1_valid),
    .io_CarryDepenIn_1_bits_taskID(Loop_1_io_CarryDepenIn_1_bits_taskID),
    .io_CarryDepenIn_1_bits_data(Loop_1_io_CarryDepenIn_1_bits_data),
    .io_CarryDepenOut_field1_0_ready(Loop_1_io_CarryDepenOut_field1_0_ready),
    .io_CarryDepenOut_field1_0_valid(Loop_1_io_CarryDepenOut_field1_0_valid),
    .io_CarryDepenOut_field1_0_bits_taskID(Loop_1_io_CarryDepenOut_field1_0_bits_taskID),
    .io_CarryDepenOut_field1_0_bits_data(Loop_1_io_CarryDepenOut_field1_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_1_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_1_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_1_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_1_io_CarryDepenOut_field0_0_bits_data),
    .io_InLiveOut_0_ready(Loop_1_io_InLiveOut_0_ready),
    .io_InLiveOut_0_valid(Loop_1_io_InLiveOut_0_valid),
    .io_InLiveOut_0_bits_taskID(Loop_1_io_InLiveOut_0_bits_taskID),
    .io_InLiveOut_0_bits_data(Loop_1_io_InLiveOut_0_bits_data),
    .io_OutLiveOut_field0_0_ready(Loop_1_io_OutLiveOut_field0_0_ready),
    .io_OutLiveOut_field0_0_valid(Loop_1_io_OutLiveOut_field0_0_valid),
    .io_OutLiveOut_field0_0_bits_taskID(Loop_1_io_OutLiveOut_field0_0_bits_taskID),
    .io_OutLiveOut_field0_0_bits_data(Loop_1_io_OutLiveOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_1_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_1_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_1_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_1_io_loopExit_0_bits_control)
  );
  LoopBlockNode_2 Loop_2 ( // @[extracted_function_reduction.scala 66:22]
    .clock(Loop_2_clock),
    .reset(Loop_2_reset),
    .io_enable_ready(Loop_2_io_enable_ready),
    .io_enable_valid(Loop_2_io_enable_valid),
    .io_enable_bits_taskID(Loop_2_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_2_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_2_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_2_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_2_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_2_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_2_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_predicate(Loop_2_io_InLiveIn_1_bits_predicate),
    .io_InLiveIn_1_bits_taskID(Loop_2_io_InLiveIn_1_bits_taskID),
    .io_InLiveIn_1_bits_data(Loop_2_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_2_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_2_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_2_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_2_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_2_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_data(Loop_2_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_2_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_2_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_taskID(Loop_2_io_InLiveIn_4_bits_taskID),
    .io_InLiveIn_4_bits_data(Loop_2_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_2_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_2_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_data(Loop_2_io_InLiveIn_5_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_2_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_2_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_data(Loop_2_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_2_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_2_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_taskID(Loop_2_io_OutLiveIn_field4_0_bits_taskID),
    .io_OutLiveIn_field4_0_bits_data(Loop_2_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_2_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_2_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_data(Loop_2_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_2_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_2_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_2_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_2_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_2_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_predicate(Loop_2_io_OutLiveIn_field1_0_bits_predicate),
    .io_OutLiveIn_field1_0_bits_taskID(Loop_2_io_OutLiveIn_field1_0_bits_taskID),
    .io_OutLiveIn_field1_0_bits_data(Loop_2_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field1_1_ready(Loop_2_io_OutLiveIn_field1_1_ready),
    .io_OutLiveIn_field1_1_valid(Loop_2_io_OutLiveIn_field1_1_valid),
    .io_OutLiveIn_field1_1_bits_taskID(Loop_2_io_OutLiveIn_field1_1_bits_taskID),
    .io_OutLiveIn_field1_1_bits_data(Loop_2_io_OutLiveIn_field1_1_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_2_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_2_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_2_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_2_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_2_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_2_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_2_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_2_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_2_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_2_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_2_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_2_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_2_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_2_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_2_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_2_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_2_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_2_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_2_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_2_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_2_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_2_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_2_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_2_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_2_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_2_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_2_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_2_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_2_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_2_io_loopExit_0_bits_control)
  );
  LoopBlockNode_3 Loop_3 ( // @[extracted_function_reduction.scala 68:22]
    .clock(Loop_3_clock),
    .reset(Loop_3_reset),
    .io_enable_ready(Loop_3_io_enable_ready),
    .io_enable_valid(Loop_3_io_enable_valid),
    .io_enable_bits_taskID(Loop_3_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_3_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_3_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_3_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_3_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_3_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_3_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_3_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_3_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_3_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_3_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_3_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_3_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_data(Loop_3_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_3_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_3_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_taskID(Loop_3_io_InLiveIn_4_bits_taskID),
    .io_InLiveIn_4_bits_data(Loop_3_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_3_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_3_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_taskID(Loop_3_io_InLiveIn_5_bits_taskID),
    .io_InLiveIn_5_bits_data(Loop_3_io_InLiveIn_5_bits_data),
    .io_InLiveIn_6_ready(Loop_3_io_InLiveIn_6_ready),
    .io_InLiveIn_6_valid(Loop_3_io_InLiveIn_6_valid),
    .io_InLiveIn_6_bits_data(Loop_3_io_InLiveIn_6_bits_data),
    .io_InLiveIn_7_ready(Loop_3_io_InLiveIn_7_ready),
    .io_InLiveIn_7_valid(Loop_3_io_InLiveIn_7_valid),
    .io_InLiveIn_7_bits_data(Loop_3_io_InLiveIn_7_bits_data),
    .io_InLiveIn_8_ready(Loop_3_io_InLiveIn_8_ready),
    .io_InLiveIn_8_valid(Loop_3_io_InLiveIn_8_valid),
    .io_InLiveIn_8_bits_taskID(Loop_3_io_InLiveIn_8_bits_taskID),
    .io_InLiveIn_8_bits_data(Loop_3_io_InLiveIn_8_bits_data),
    .io_OutLiveIn_field8_0_ready(Loop_3_io_OutLiveIn_field8_0_ready),
    .io_OutLiveIn_field8_0_valid(Loop_3_io_OutLiveIn_field8_0_valid),
    .io_OutLiveIn_field8_0_bits_taskID(Loop_3_io_OutLiveIn_field8_0_bits_taskID),
    .io_OutLiveIn_field8_0_bits_data(Loop_3_io_OutLiveIn_field8_0_bits_data),
    .io_OutLiveIn_field8_1_ready(Loop_3_io_OutLiveIn_field8_1_ready),
    .io_OutLiveIn_field8_1_valid(Loop_3_io_OutLiveIn_field8_1_valid),
    .io_OutLiveIn_field8_1_bits_data(Loop_3_io_OutLiveIn_field8_1_bits_data),
    .io_OutLiveIn_field7_0_ready(Loop_3_io_OutLiveIn_field7_0_ready),
    .io_OutLiveIn_field7_0_valid(Loop_3_io_OutLiveIn_field7_0_valid),
    .io_OutLiveIn_field7_0_bits_data(Loop_3_io_OutLiveIn_field7_0_bits_data),
    .io_OutLiveIn_field6_0_ready(Loop_3_io_OutLiveIn_field6_0_ready),
    .io_OutLiveIn_field6_0_valid(Loop_3_io_OutLiveIn_field6_0_valid),
    .io_OutLiveIn_field6_0_bits_data(Loop_3_io_OutLiveIn_field6_0_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_3_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_3_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_taskID(Loop_3_io_OutLiveIn_field5_0_bits_taskID),
    .io_OutLiveIn_field5_0_bits_data(Loop_3_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_3_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_3_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_taskID(Loop_3_io_OutLiveIn_field4_0_bits_taskID),
    .io_OutLiveIn_field4_0_bits_data(Loop_3_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_3_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_3_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_data(Loop_3_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_3_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_3_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_3_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_3_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_3_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_3_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_3_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_3_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_3_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_3_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_3_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_3_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_3_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_3_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_3_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_3_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_3_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_3_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_3_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_3_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_3_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_3_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_3_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_3_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_3_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_3_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_3_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_3_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_3_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_3_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_3_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_3_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_3_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_3_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_3_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_3_io_loopExit_0_bits_control)
  );
  LoopBlockNode_4 Loop_4 ( // @[extracted_function_reduction.scala 70:22]
    .clock(Loop_4_clock),
    .reset(Loop_4_reset),
    .io_enable_ready(Loop_4_io_enable_ready),
    .io_enable_valid(Loop_4_io_enable_valid),
    .io_enable_bits_taskID(Loop_4_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_4_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_4_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_4_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_4_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_4_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_4_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_4_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_4_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_4_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_4_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_4_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_4_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_taskID(Loop_4_io_InLiveIn_3_bits_taskID),
    .io_InLiveIn_3_bits_data(Loop_4_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_4_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_4_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_taskID(Loop_4_io_InLiveIn_4_bits_taskID),
    .io_InLiveIn_4_bits_data(Loop_4_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_4_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_4_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_data(Loop_4_io_InLiveIn_5_bits_data),
    .io_InLiveIn_6_ready(Loop_4_io_InLiveIn_6_ready),
    .io_InLiveIn_6_valid(Loop_4_io_InLiveIn_6_valid),
    .io_InLiveIn_6_bits_data(Loop_4_io_InLiveIn_6_bits_data),
    .io_InLiveIn_7_ready(Loop_4_io_InLiveIn_7_ready),
    .io_InLiveIn_7_valid(Loop_4_io_InLiveIn_7_valid),
    .io_InLiveIn_7_bits_taskID(Loop_4_io_InLiveIn_7_bits_taskID),
    .io_InLiveIn_7_bits_data(Loop_4_io_InLiveIn_7_bits_data),
    .io_InLiveIn_8_ready(Loop_4_io_InLiveIn_8_ready),
    .io_InLiveIn_8_valid(Loop_4_io_InLiveIn_8_valid),
    .io_InLiveIn_8_bits_taskID(Loop_4_io_InLiveIn_8_bits_taskID),
    .io_InLiveIn_8_bits_data(Loop_4_io_InLiveIn_8_bits_data),
    .io_InLiveIn_9_ready(Loop_4_io_InLiveIn_9_ready),
    .io_InLiveIn_9_valid(Loop_4_io_InLiveIn_9_valid),
    .io_InLiveIn_9_bits_data(Loop_4_io_InLiveIn_9_bits_data),
    .io_InLiveIn_10_ready(Loop_4_io_InLiveIn_10_ready),
    .io_InLiveIn_10_valid(Loop_4_io_InLiveIn_10_valid),
    .io_InLiveIn_10_bits_taskID(Loop_4_io_InLiveIn_10_bits_taskID),
    .io_InLiveIn_10_bits_data(Loop_4_io_InLiveIn_10_bits_data),
    .io_InLiveIn_11_ready(Loop_4_io_InLiveIn_11_ready),
    .io_InLiveIn_11_valid(Loop_4_io_InLiveIn_11_valid),
    .io_InLiveIn_11_bits_data(Loop_4_io_InLiveIn_11_bits_data),
    .io_OutLiveIn_field11_0_ready(Loop_4_io_OutLiveIn_field11_0_ready),
    .io_OutLiveIn_field11_0_valid(Loop_4_io_OutLiveIn_field11_0_valid),
    .io_OutLiveIn_field11_0_bits_data(Loop_4_io_OutLiveIn_field11_0_bits_data),
    .io_OutLiveIn_field10_0_ready(Loop_4_io_OutLiveIn_field10_0_ready),
    .io_OutLiveIn_field10_0_valid(Loop_4_io_OutLiveIn_field10_0_valid),
    .io_OutLiveIn_field10_0_bits_taskID(Loop_4_io_OutLiveIn_field10_0_bits_taskID),
    .io_OutLiveIn_field10_0_bits_data(Loop_4_io_OutLiveIn_field10_0_bits_data),
    .io_OutLiveIn_field10_1_ready(Loop_4_io_OutLiveIn_field10_1_ready),
    .io_OutLiveIn_field10_1_valid(Loop_4_io_OutLiveIn_field10_1_valid),
    .io_OutLiveIn_field10_1_bits_data(Loop_4_io_OutLiveIn_field10_1_bits_data),
    .io_OutLiveIn_field9_0_ready(Loop_4_io_OutLiveIn_field9_0_ready),
    .io_OutLiveIn_field9_0_valid(Loop_4_io_OutLiveIn_field9_0_valid),
    .io_OutLiveIn_field9_0_bits_data(Loop_4_io_OutLiveIn_field9_0_bits_data),
    .io_OutLiveIn_field8_0_ready(Loop_4_io_OutLiveIn_field8_0_ready),
    .io_OutLiveIn_field8_0_valid(Loop_4_io_OutLiveIn_field8_0_valid),
    .io_OutLiveIn_field8_0_bits_taskID(Loop_4_io_OutLiveIn_field8_0_bits_taskID),
    .io_OutLiveIn_field8_0_bits_data(Loop_4_io_OutLiveIn_field8_0_bits_data),
    .io_OutLiveIn_field7_0_ready(Loop_4_io_OutLiveIn_field7_0_ready),
    .io_OutLiveIn_field7_0_valid(Loop_4_io_OutLiveIn_field7_0_valid),
    .io_OutLiveIn_field7_0_bits_taskID(Loop_4_io_OutLiveIn_field7_0_bits_taskID),
    .io_OutLiveIn_field7_0_bits_data(Loop_4_io_OutLiveIn_field7_0_bits_data),
    .io_OutLiveIn_field6_0_ready(Loop_4_io_OutLiveIn_field6_0_ready),
    .io_OutLiveIn_field6_0_valid(Loop_4_io_OutLiveIn_field6_0_valid),
    .io_OutLiveIn_field6_0_bits_data(Loop_4_io_OutLiveIn_field6_0_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_4_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_4_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_data(Loop_4_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_4_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_4_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_taskID(Loop_4_io_OutLiveIn_field4_0_bits_taskID),
    .io_OutLiveIn_field4_0_bits_data(Loop_4_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_4_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_4_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_taskID(Loop_4_io_OutLiveIn_field3_0_bits_taskID),
    .io_OutLiveIn_field3_0_bits_data(Loop_4_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_4_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_4_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_4_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_4_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_4_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_4_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_4_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_4_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_4_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_4_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_4_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_4_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_4_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_4_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_4_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_4_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_4_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_4_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_4_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_4_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_4_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_4_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_4_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_4_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_4_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_4_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_4_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_4_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_4_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_4_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_4_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_4_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_4_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_4_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_4_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_4_io_loopExit_0_bits_control)
  );
  LoopBlockNode_5 Loop_5 ( // @[extracted_function_reduction.scala 72:22]
    .clock(Loop_5_clock),
    .reset(Loop_5_reset),
    .io_enable_ready(Loop_5_io_enable_ready),
    .io_enable_valid(Loop_5_io_enable_valid),
    .io_enable_bits_taskID(Loop_5_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_5_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_5_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_5_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_taskID(Loop_5_io_InLiveIn_0_bits_taskID),
    .io_InLiveIn_0_bits_data(Loop_5_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_5_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_5_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_5_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_5_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_5_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_taskID(Loop_5_io_InLiveIn_2_bits_taskID),
    .io_InLiveIn_2_bits_data(Loop_5_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_5_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_5_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_taskID(Loop_5_io_InLiveIn_3_bits_taskID),
    .io_InLiveIn_3_bits_data(Loop_5_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_5_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_5_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_taskID(Loop_5_io_InLiveIn_4_bits_taskID),
    .io_InLiveIn_4_bits_data(Loop_5_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_5_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_5_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_data(Loop_5_io_InLiveIn_5_bits_data),
    .io_InLiveIn_6_ready(Loop_5_io_InLiveIn_6_ready),
    .io_InLiveIn_6_valid(Loop_5_io_InLiveIn_6_valid),
    .io_InLiveIn_6_bits_taskID(Loop_5_io_InLiveIn_6_bits_taskID),
    .io_InLiveIn_6_bits_data(Loop_5_io_InLiveIn_6_bits_data),
    .io_InLiveIn_7_ready(Loop_5_io_InLiveIn_7_ready),
    .io_InLiveIn_7_valid(Loop_5_io_InLiveIn_7_valid),
    .io_InLiveIn_7_bits_data(Loop_5_io_InLiveIn_7_bits_data),
    .io_InLiveIn_8_ready(Loop_5_io_InLiveIn_8_ready),
    .io_InLiveIn_8_valid(Loop_5_io_InLiveIn_8_valid),
    .io_InLiveIn_8_bits_taskID(Loop_5_io_InLiveIn_8_bits_taskID),
    .io_InLiveIn_8_bits_data(Loop_5_io_InLiveIn_8_bits_data),
    .io_InLiveIn_9_ready(Loop_5_io_InLiveIn_9_ready),
    .io_InLiveIn_9_valid(Loop_5_io_InLiveIn_9_valid),
    .io_InLiveIn_9_bits_data(Loop_5_io_InLiveIn_9_bits_data),
    .io_InLiveIn_10_ready(Loop_5_io_InLiveIn_10_ready),
    .io_InLiveIn_10_valid(Loop_5_io_InLiveIn_10_valid),
    .io_InLiveIn_10_bits_data(Loop_5_io_InLiveIn_10_bits_data),
    .io_InLiveIn_11_ready(Loop_5_io_InLiveIn_11_ready),
    .io_InLiveIn_11_valid(Loop_5_io_InLiveIn_11_valid),
    .io_InLiveIn_11_bits_taskID(Loop_5_io_InLiveIn_11_bits_taskID),
    .io_InLiveIn_11_bits_data(Loop_5_io_InLiveIn_11_bits_data),
    .io_InLiveIn_12_ready(Loop_5_io_InLiveIn_12_ready),
    .io_InLiveIn_12_valid(Loop_5_io_InLiveIn_12_valid),
    .io_InLiveIn_12_bits_data(Loop_5_io_InLiveIn_12_bits_data),
    .io_InLiveIn_13_ready(Loop_5_io_InLiveIn_13_ready),
    .io_InLiveIn_13_valid(Loop_5_io_InLiveIn_13_valid),
    .io_InLiveIn_13_bits_data(Loop_5_io_InLiveIn_13_bits_data),
    .io_InLiveIn_14_ready(Loop_5_io_InLiveIn_14_ready),
    .io_InLiveIn_14_valid(Loop_5_io_InLiveIn_14_valid),
    .io_InLiveIn_14_bits_data(Loop_5_io_InLiveIn_14_bits_data),
    .io_OutLiveIn_field14_0_ready(Loop_5_io_OutLiveIn_field14_0_ready),
    .io_OutLiveIn_field14_0_valid(Loop_5_io_OutLiveIn_field14_0_valid),
    .io_OutLiveIn_field14_0_bits_data(Loop_5_io_OutLiveIn_field14_0_bits_data),
    .io_OutLiveIn_field13_0_ready(Loop_5_io_OutLiveIn_field13_0_ready),
    .io_OutLiveIn_field13_0_valid(Loop_5_io_OutLiveIn_field13_0_valid),
    .io_OutLiveIn_field13_0_bits_data(Loop_5_io_OutLiveIn_field13_0_bits_data),
    .io_OutLiveIn_field12_0_ready(Loop_5_io_OutLiveIn_field12_0_ready),
    .io_OutLiveIn_field12_0_valid(Loop_5_io_OutLiveIn_field12_0_valid),
    .io_OutLiveIn_field12_0_bits_data(Loop_5_io_OutLiveIn_field12_0_bits_data),
    .io_OutLiveIn_field11_0_ready(Loop_5_io_OutLiveIn_field11_0_ready),
    .io_OutLiveIn_field11_0_valid(Loop_5_io_OutLiveIn_field11_0_valid),
    .io_OutLiveIn_field11_0_bits_taskID(Loop_5_io_OutLiveIn_field11_0_bits_taskID),
    .io_OutLiveIn_field11_0_bits_data(Loop_5_io_OutLiveIn_field11_0_bits_data),
    .io_OutLiveIn_field10_0_ready(Loop_5_io_OutLiveIn_field10_0_ready),
    .io_OutLiveIn_field10_0_valid(Loop_5_io_OutLiveIn_field10_0_valid),
    .io_OutLiveIn_field10_0_bits_data(Loop_5_io_OutLiveIn_field10_0_bits_data),
    .io_OutLiveIn_field9_0_ready(Loop_5_io_OutLiveIn_field9_0_ready),
    .io_OutLiveIn_field9_0_valid(Loop_5_io_OutLiveIn_field9_0_valid),
    .io_OutLiveIn_field9_0_bits_data(Loop_5_io_OutLiveIn_field9_0_bits_data),
    .io_OutLiveIn_field8_0_ready(Loop_5_io_OutLiveIn_field8_0_ready),
    .io_OutLiveIn_field8_0_valid(Loop_5_io_OutLiveIn_field8_0_valid),
    .io_OutLiveIn_field8_0_bits_taskID(Loop_5_io_OutLiveIn_field8_0_bits_taskID),
    .io_OutLiveIn_field8_0_bits_data(Loop_5_io_OutLiveIn_field8_0_bits_data),
    .io_OutLiveIn_field7_0_ready(Loop_5_io_OutLiveIn_field7_0_ready),
    .io_OutLiveIn_field7_0_valid(Loop_5_io_OutLiveIn_field7_0_valid),
    .io_OutLiveIn_field7_0_bits_data(Loop_5_io_OutLiveIn_field7_0_bits_data),
    .io_OutLiveIn_field6_0_ready(Loop_5_io_OutLiveIn_field6_0_ready),
    .io_OutLiveIn_field6_0_valid(Loop_5_io_OutLiveIn_field6_0_valid),
    .io_OutLiveIn_field6_0_bits_taskID(Loop_5_io_OutLiveIn_field6_0_bits_taskID),
    .io_OutLiveIn_field6_0_bits_data(Loop_5_io_OutLiveIn_field6_0_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_5_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_5_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_data(Loop_5_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_5_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_5_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_taskID(Loop_5_io_OutLiveIn_field4_0_bits_taskID),
    .io_OutLiveIn_field4_0_bits_data(Loop_5_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_5_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_5_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_taskID(Loop_5_io_OutLiveIn_field3_0_bits_taskID),
    .io_OutLiveIn_field3_0_bits_data(Loop_5_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_5_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_5_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_taskID(Loop_5_io_OutLiveIn_field2_0_bits_taskID),
    .io_OutLiveIn_field2_0_bits_data(Loop_5_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_5_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_5_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_5_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_5_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_5_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_taskID(Loop_5_io_OutLiveIn_field0_0_bits_taskID),
    .io_OutLiveIn_field0_0_bits_data(Loop_5_io_OutLiveIn_field0_0_bits_data),
    .io_OutLiveIn_field0_1_ready(Loop_5_io_OutLiveIn_field0_1_ready),
    .io_OutLiveIn_field0_1_valid(Loop_5_io_OutLiveIn_field0_1_valid),
    .io_OutLiveIn_field0_1_bits_data(Loop_5_io_OutLiveIn_field0_1_bits_data),
    .io_activate_loop_start_ready(Loop_5_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_5_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_5_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_5_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_5_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_5_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_5_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_5_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_5_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_5_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_5_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_5_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_5_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_5_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_5_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_5_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_5_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_5_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_5_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_5_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_5_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_5_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_5_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_5_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_5_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_5_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_5_io_loopExit_0_bits_control)
  );
  BasicBlockNoMaskFastNode bb_entry0 ( // @[extracted_function_reduction.scala 80:25]
    .clock(bb_entry0_clock),
    .reset(bb_entry0_reset),
    .io_predicateIn_0_ready(bb_entry0_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_entry0_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_entry0_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_entry0_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_entry0_io_Out_0_ready),
    .io_Out_0_valid(bb_entry0_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_entry0_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_entry0_io_Out_0_bits_control),
    .io_Out_1_ready(bb_entry0_io_Out_1_ready),
    .io_Out_1_valid(bb_entry0_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_entry0_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_entry0_io_Out_1_bits_control),
    .io_Out_2_ready(bb_entry0_io_Out_2_ready),
    .io_Out_2_valid(bb_entry0_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_entry0_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_entry0_io_Out_2_bits_control)
  );
  BasicBlockNoMaskFastNode_1 bb_for_body_lr_ph1 ( // @[extracted_function_reduction.scala 82:34]
    .clock(bb_for_body_lr_ph1_clock),
    .reset(bb_for_body_lr_ph1_reset),
    .io_predicateIn_0_ready(bb_for_body_lr_ph1_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body_lr_ph1_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body_lr_ph1_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body_lr_ph1_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_body_lr_ph1_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body_lr_ph1_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body_lr_ph1_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_body_lr_ph1_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_body_lr_ph1_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body_lr_ph1_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body_lr_ph1_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_body_lr_ph1_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_body_lr_ph1_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body_lr_ph1_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body_lr_ph1_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_body_lr_ph1_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_body_lr_ph1_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body_lr_ph1_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_body_lr_ph1_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_body_lr_ph1_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_body_lr_ph1_io_Out_4_ready),
    .io_Out_4_valid(bb_for_body_lr_ph1_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_body_lr_ph1_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_body_lr_ph1_io_Out_4_bits_control)
  );
  BasicBlockNoMaskFastNode_2 bb_for_cond_cleanup_loopexit2 ( // @[extracted_function_reduction.scala 84:45]
    .clock(bb_for_cond_cleanup_loopexit2_clock),
    .reset(bb_for_cond_cleanup_loopexit2_reset),
    .io_predicateIn_0_ready(bb_for_cond_cleanup_loopexit2_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup_loopexit2_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup_loopexit2_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup_loopexit2_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_cond_cleanup_loopexit2_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup_loopexit2_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup_loopexit2_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_cond_cleanup_loopexit2_io_Out_0_bits_control)
  );
  BasicBlockNoMaskFastNode_3 bb_for_cond_cleanup3 ( // @[extracted_function_reduction.scala 86:36]
    .clock(bb_for_cond_cleanup3_clock),
    .reset(bb_for_cond_cleanup3_reset),
    .io_predicateIn_0_ready(bb_for_cond_cleanup3_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup3_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup3_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup3_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_cond_cleanup3_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_cond_cleanup3_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_cond_cleanup3_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_cond_cleanup3_io_predicateIn_1_bits_control),
    .io_Out_0_ready(bb_for_cond_cleanup3_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup3_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup3_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_cond_cleanup3_io_Out_0_bits_control)
  );
  BasicBlockNode bb_for_body4 ( // @[extracted_function_reduction.scala 88:28]
    .clock(bb_for_body4_clock),
    .reset(bb_for_body4_reset),
    .io_MaskBB_0_ready(bb_for_body4_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body4_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body4_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_for_body4_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body4_io_Out_0_valid),
    .io_Out_0_bits_control(bb_for_body4_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_body4_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body4_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body4_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_body4_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_body4_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body4_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body4_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_body4_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_body4_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body4_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_body4_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_body4_io_Out_3_bits_control),
    .io_predicateIn_0_ready(bb_for_body4_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body4_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body4_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body4_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body4_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body4_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body4_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body4_io_predicateIn_1_bits_control)
  );
  BasicBlockNoMaskFastNode_4 bb_for_body7_preheader5 ( // @[extracted_function_reduction.scala 90:39]
    .clock(bb_for_body7_preheader5_clock),
    .reset(bb_for_body7_preheader5_reset),
    .io_predicateIn_0_ready(bb_for_body7_preheader5_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body7_preheader5_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body7_preheader5_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body7_preheader5_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_body7_preheader5_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body7_preheader5_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body7_preheader5_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_body7_preheader5_io_Out_0_bits_control)
  );
  BasicBlockNoMaskFastNode_5 bb_for_cond_cleanup6_loopexit6 ( // @[extracted_function_reduction.scala 92:46]
    .clock(bb_for_cond_cleanup6_loopexit6_clock),
    .reset(bb_for_cond_cleanup6_loopexit6_reset),
    .io_predicateIn_0_ready(bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_cond_cleanup6_loopexit6_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup6_loopexit6_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup6_loopexit6_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_cond_cleanup6_loopexit6_io_Out_0_bits_control)
  );
  BasicBlockNoMaskFastNode_6 bb_for_cond_cleanup67 ( // @[extracted_function_reduction.scala 94:37]
    .clock(bb_for_cond_cleanup67_clock),
    .reset(bb_for_cond_cleanup67_reset),
    .io_predicateIn_0_ready(bb_for_cond_cleanup67_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup67_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup67_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup67_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_cond_cleanup67_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_cond_cleanup67_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_cond_cleanup67_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_cond_cleanup67_io_predicateIn_1_bits_control),
    .io_Out_0_ready(bb_for_cond_cleanup67_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup67_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup67_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_cond_cleanup67_io_Out_1_ready),
    .io_Out_1_valid(bb_for_cond_cleanup67_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_cond_cleanup67_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_cond_cleanup67_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_cond_cleanup67_io_Out_2_ready),
    .io_Out_2_valid(bb_for_cond_cleanup67_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_cond_cleanup67_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_cond_cleanup67_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_cond_cleanup67_io_Out_3_ready),
    .io_Out_3_valid(bb_for_cond_cleanup67_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_cond_cleanup67_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_cond_cleanup67_io_Out_3_bits_control)
  );
  BasicBlockNode_1 bb_for_body78 ( // @[extracted_function_reduction.scala 96:29]
    .clock(bb_for_body78_clock),
    .reset(bb_for_body78_reset),
    .io_MaskBB_0_ready(bb_for_body78_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body78_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body78_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_for_body78_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body78_io_Out_0_valid),
    .io_Out_0_bits_control(bb_for_body78_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_body78_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body78_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body78_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_body78_io_Out_1_bits_control),
    .io_predicateIn_0_ready(bb_for_body78_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body78_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body78_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body78_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body78_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body78_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body78_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body78_io_predicateIn_1_bits_control)
  );
  BasicBlockNoMaskFastNode_7 bb_for_body15_lr_ph9 ( // @[extracted_function_reduction.scala 98:36]
    .clock(bb_for_body15_lr_ph9_clock),
    .reset(bb_for_body15_lr_ph9_reset),
    .io_predicateIn_0_ready(bb_for_body15_lr_ph9_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body15_lr_ph9_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body15_lr_ph9_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body15_lr_ph9_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_body15_lr_ph9_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body15_lr_ph9_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body15_lr_ph9_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_body15_lr_ph9_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_body15_lr_ph9_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body15_lr_ph9_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body15_lr_ph9_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_body15_lr_ph9_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_body15_lr_ph9_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body15_lr_ph9_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body15_lr_ph9_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_body15_lr_ph9_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_body15_lr_ph9_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body15_lr_ph9_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_body15_lr_ph9_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_body15_lr_ph9_io_Out_3_bits_control)
  );
  BasicBlockNoMaskFastNode_8 bb_for_cond_cleanup14_loopexit10 ( // @[extracted_function_reduction.scala 100:48]
    .clock(bb_for_cond_cleanup14_loopexit10_clock),
    .reset(bb_for_cond_cleanup14_loopexit10_reset),
    .io_predicateIn_0_ready(bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_cond_cleanup14_loopexit10_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup14_loopexit10_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup14_loopexit10_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_cond_cleanup14_loopexit10_io_Out_0_bits_control)
  );
  BasicBlockNoMaskFastNode_9 bb_for_cond_cleanup1411 ( // @[extracted_function_reduction.scala 102:39]
    .clock(bb_for_cond_cleanup1411_clock),
    .reset(bb_for_cond_cleanup1411_reset),
    .io_predicateIn_0_ready(bb_for_cond_cleanup1411_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup1411_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup1411_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup1411_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_cond_cleanup1411_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_cond_cleanup1411_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_cond_cleanup1411_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_cond_cleanup1411_io_predicateIn_1_bits_control),
    .io_Out_0_ready(bb_for_cond_cleanup1411_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup1411_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup1411_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_cond_cleanup1411_io_Out_1_ready),
    .io_Out_1_valid(bb_for_cond_cleanup1411_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_cond_cleanup1411_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_cond_cleanup1411_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_cond_cleanup1411_io_Out_2_ready),
    .io_Out_2_valid(bb_for_cond_cleanup1411_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_cond_cleanup1411_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_cond_cleanup1411_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_cond_cleanup1411_io_Out_3_ready),
    .io_Out_3_valid(bb_for_cond_cleanup1411_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_cond_cleanup1411_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_cond_cleanup1411_io_Out_3_bits_control)
  );
  BasicBlockNode_2 bb_for_body1512 ( // @[extracted_function_reduction.scala 104:31]
    .clock(bb_for_body1512_clock),
    .reset(bb_for_body1512_reset),
    .io_MaskBB_0_ready(bb_for_body1512_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body1512_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body1512_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_for_body1512_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body1512_io_Out_0_valid),
    .io_Out_0_bits_control(bb_for_body1512_io_Out_0_bits_control),
    .io_Out_1_ready(bb_for_body1512_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body1512_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body1512_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_body1512_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_body1512_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body1512_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body1512_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_body1512_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_body1512_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body1512_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_body1512_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_body1512_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_body1512_io_Out_4_ready),
    .io_Out_4_valid(bb_for_body1512_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_body1512_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_body1512_io_Out_4_bits_control),
    .io_Out_5_ready(bb_for_body1512_io_Out_5_ready),
    .io_Out_5_valid(bb_for_body1512_io_Out_5_valid),
    .io_Out_5_bits_taskID(bb_for_body1512_io_Out_5_bits_taskID),
    .io_Out_5_bits_control(bb_for_body1512_io_Out_5_bits_control),
    .io_predicateIn_0_ready(bb_for_body1512_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body1512_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body1512_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body1512_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body1512_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body1512_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body1512_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body1512_io_predicateIn_1_bits_control)
  );
  BasicBlockNoMaskFastNode_10 bb_for_cond_cleanup2013 ( // @[extracted_function_reduction.scala 106:39]
    .clock(bb_for_cond_cleanup2013_clock),
    .reset(bb_for_cond_cleanup2013_reset),
    .io_predicateIn_0_ready(bb_for_cond_cleanup2013_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup2013_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup2013_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup2013_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_cond_cleanup2013_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup2013_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup2013_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_cond_cleanup2013_io_Out_1_ready),
    .io_Out_1_valid(bb_for_cond_cleanup2013_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_cond_cleanup2013_io_Out_1_bits_taskID),
    .io_Out_1_bits_control(bb_for_cond_cleanup2013_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_cond_cleanup2013_io_Out_2_ready),
    .io_Out_2_valid(bb_for_cond_cleanup2013_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_cond_cleanup2013_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_cond_cleanup2013_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_cond_cleanup2013_io_Out_3_ready),
    .io_Out_3_valid(bb_for_cond_cleanup2013_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_cond_cleanup2013_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_cond_cleanup2013_io_Out_3_bits_control)
  );
  BasicBlockNode_3 bb_for_body2114 ( // @[extracted_function_reduction.scala 108:31]
    .clock(bb_for_body2114_clock),
    .reset(bb_for_body2114_reset),
    .io_MaskBB_0_ready(bb_for_body2114_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body2114_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body2114_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_for_body2114_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body2114_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body2114_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_body2114_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body2114_io_Out_1_valid),
    .io_Out_1_bits_control(bb_for_body2114_io_Out_1_bits_control),
    .io_Out_2_ready(bb_for_body2114_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body2114_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body2114_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_body2114_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_body2114_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body2114_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_body2114_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_body2114_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_body2114_io_Out_4_ready),
    .io_Out_4_valid(bb_for_body2114_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_body2114_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_body2114_io_Out_4_bits_control),
    .io_predicateIn_0_ready(bb_for_body2114_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body2114_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body2114_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body2114_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body2114_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body2114_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body2114_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body2114_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_4 bb_for_cond_cleanup2615 ( // @[extracted_function_reduction.scala 110:39]
    .clock(bb_for_cond_cleanup2615_clock),
    .reset(bb_for_cond_cleanup2615_reset),
    .io_Out_0_ready(bb_for_cond_cleanup2615_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup2615_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup2615_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_cond_cleanup2615_io_Out_1_ready),
    .io_Out_1_valid(bb_for_cond_cleanup2615_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_cond_cleanup2615_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_for_cond_cleanup2615_io_Out_2_ready),
    .io_Out_2_valid(bb_for_cond_cleanup2615_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_cond_cleanup2615_io_Out_2_bits_taskID),
    .io_Out_3_ready(bb_for_cond_cleanup2615_io_Out_3_ready),
    .io_Out_3_valid(bb_for_cond_cleanup2615_io_Out_3_valid),
    .io_Out_3_bits_control(bb_for_cond_cleanup2615_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_cond_cleanup2615_io_Out_4_ready),
    .io_Out_4_valid(bb_for_cond_cleanup2615_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_cond_cleanup2615_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_cond_cleanup2615_io_Out_4_bits_control),
    .io_Out_5_ready(bb_for_cond_cleanup2615_io_Out_5_ready),
    .io_Out_5_valid(bb_for_cond_cleanup2615_io_Out_5_valid),
    .io_Out_5_bits_taskID(bb_for_cond_cleanup2615_io_Out_5_bits_taskID),
    .io_Out_6_ready(bb_for_cond_cleanup2615_io_Out_6_ready),
    .io_Out_6_valid(bb_for_cond_cleanup2615_io_Out_6_valid),
    .io_Out_6_bits_taskID(bb_for_cond_cleanup2615_io_Out_6_bits_taskID),
    .io_Out_6_bits_control(bb_for_cond_cleanup2615_io_Out_6_bits_control),
    .io_Out_7_ready(bb_for_cond_cleanup2615_io_Out_7_ready),
    .io_Out_7_valid(bb_for_cond_cleanup2615_io_Out_7_valid),
    .io_Out_7_bits_taskID(bb_for_cond_cleanup2615_io_Out_7_bits_taskID),
    .io_Out_7_bits_control(bb_for_cond_cleanup2615_io_Out_7_bits_control),
    .io_Out_8_ready(bb_for_cond_cleanup2615_io_Out_8_ready),
    .io_Out_8_valid(bb_for_cond_cleanup2615_io_Out_8_valid),
    .io_Out_8_bits_taskID(bb_for_cond_cleanup2615_io_Out_8_bits_taskID),
    .io_Out_8_bits_control(bb_for_cond_cleanup2615_io_Out_8_bits_control),
    .io_Out_9_ready(bb_for_cond_cleanup2615_io_Out_9_ready),
    .io_Out_9_valid(bb_for_cond_cleanup2615_io_Out_9_valid),
    .io_Out_9_bits_taskID(bb_for_cond_cleanup2615_io_Out_9_bits_taskID),
    .io_Out_9_bits_control(bb_for_cond_cleanup2615_io_Out_9_bits_control),
    .io_Out_10_ready(bb_for_cond_cleanup2615_io_Out_10_ready),
    .io_Out_10_valid(bb_for_cond_cleanup2615_io_Out_10_valid),
    .io_Out_10_bits_taskID(bb_for_cond_cleanup2615_io_Out_10_bits_taskID),
    .io_Out_10_bits_control(bb_for_cond_cleanup2615_io_Out_10_bits_control),
    .io_Out_11_ready(bb_for_cond_cleanup2615_io_Out_11_ready),
    .io_Out_11_valid(bb_for_cond_cleanup2615_io_Out_11_valid),
    .io_Out_11_bits_taskID(bb_for_cond_cleanup2615_io_Out_11_bits_taskID),
    .io_Out_11_bits_control(bb_for_cond_cleanup2615_io_Out_11_bits_control),
    .io_predicateIn_0_ready(bb_for_cond_cleanup2615_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup2615_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup2615_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup2615_io_predicateIn_0_bits_control)
  );
  BasicBlockNode_5 bb_for_body2716 ( // @[extracted_function_reduction.scala 112:31]
    .clock(bb_for_body2716_clock),
    .reset(bb_for_body2716_reset),
    .io_MaskBB_0_ready(bb_for_body2716_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body2716_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body2716_io_MaskBB_0_bits),
    .io_MaskBB_1_ready(bb_for_body2716_io_MaskBB_1_ready),
    .io_MaskBB_1_valid(bb_for_body2716_io_MaskBB_1_valid),
    .io_MaskBB_1_bits(bb_for_body2716_io_MaskBB_1_bits),
    .io_Out_0_ready(bb_for_body2716_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body2716_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body2716_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_body2716_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body2716_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body2716_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_for_body2716_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body2716_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body2716_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_body2716_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_body2716_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body2716_io_Out_3_valid),
    .io_Out_3_bits_control(bb_for_body2716_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_body2716_io_Out_4_ready),
    .io_Out_4_valid(bb_for_body2716_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_body2716_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_body2716_io_Out_4_bits_control),
    .io_Out_5_ready(bb_for_body2716_io_Out_5_ready),
    .io_Out_5_valid(bb_for_body2716_io_Out_5_valid),
    .io_Out_5_bits_taskID(bb_for_body2716_io_Out_5_bits_taskID),
    .io_Out_5_bits_control(bb_for_body2716_io_Out_5_bits_control),
    .io_Out_6_ready(bb_for_body2716_io_Out_6_ready),
    .io_Out_6_valid(bb_for_body2716_io_Out_6_valid),
    .io_Out_6_bits_taskID(bb_for_body2716_io_Out_6_bits_taskID),
    .io_Out_6_bits_control(bb_for_body2716_io_Out_6_bits_control),
    .io_Out_7_ready(bb_for_body2716_io_Out_7_ready),
    .io_Out_7_valid(bb_for_body2716_io_Out_7_valid),
    .io_Out_7_bits_taskID(bb_for_body2716_io_Out_7_bits_taskID),
    .io_Out_7_bits_control(bb_for_body2716_io_Out_7_bits_control),
    .io_predicateIn_0_ready(bb_for_body2716_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body2716_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body2716_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body2716_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body2716_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body2716_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body2716_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body2716_io_predicateIn_1_bits_control)
  );
  BasicBlockNode_6 bb_for_cond_cleanup3317 ( // @[extracted_function_reduction.scala 114:39]
    .clock(bb_for_cond_cleanup3317_clock),
    .reset(bb_for_cond_cleanup3317_reset),
    .io_Out_0_ready(bb_for_cond_cleanup3317_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup3317_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup3317_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_cond_cleanup3317_io_Out_1_ready),
    .io_Out_1_valid(bb_for_cond_cleanup3317_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_cond_cleanup3317_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_for_cond_cleanup3317_io_Out_2_ready),
    .io_Out_2_valid(bb_for_cond_cleanup3317_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_cond_cleanup3317_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_cond_cleanup3317_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_cond_cleanup3317_io_Out_3_ready),
    .io_Out_3_valid(bb_for_cond_cleanup3317_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_cond_cleanup3317_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_cond_cleanup3317_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_cond_cleanup3317_io_Out_4_ready),
    .io_Out_4_valid(bb_for_cond_cleanup3317_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_cond_cleanup3317_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_cond_cleanup3317_io_Out_4_bits_control),
    .io_Out_5_ready(bb_for_cond_cleanup3317_io_Out_5_ready),
    .io_Out_5_valid(bb_for_cond_cleanup3317_io_Out_5_valid),
    .io_Out_5_bits_taskID(bb_for_cond_cleanup3317_io_Out_5_bits_taskID),
    .io_Out_5_bits_control(bb_for_cond_cleanup3317_io_Out_5_bits_control),
    .io_predicateIn_0_ready(bb_for_cond_cleanup3317_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup3317_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup3317_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup3317_io_predicateIn_0_bits_control)
  );
  BasicBlockNode_7 bb_for_body3418 ( // @[extracted_function_reduction.scala 116:31]
    .clock(bb_for_body3418_clock),
    .reset(bb_for_body3418_reset),
    .io_MaskBB_0_ready(bb_for_body3418_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body3418_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body3418_io_MaskBB_0_bits),
    .io_MaskBB_1_ready(bb_for_body3418_io_MaskBB_1_ready),
    .io_MaskBB_1_valid(bb_for_body3418_io_MaskBB_1_valid),
    .io_MaskBB_1_bits(bb_for_body3418_io_MaskBB_1_bits),
    .io_Out_0_ready(bb_for_body3418_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body3418_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body3418_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_body3418_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body3418_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body3418_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_for_body3418_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body3418_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body3418_io_Out_2_bits_taskID),
    .io_Out_3_ready(bb_for_body3418_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body3418_io_Out_3_valid),
    .io_Out_3_bits_control(bb_for_body3418_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_body3418_io_Out_4_ready),
    .io_Out_4_valid(bb_for_body3418_io_Out_4_valid),
    .io_Out_4_bits_control(bb_for_body3418_io_Out_4_bits_control),
    .io_Out_5_ready(bb_for_body3418_io_Out_5_ready),
    .io_Out_5_valid(bb_for_body3418_io_Out_5_valid),
    .io_Out_5_bits_taskID(bb_for_body3418_io_Out_5_bits_taskID),
    .io_Out_5_bits_control(bb_for_body3418_io_Out_5_bits_control),
    .io_Out_6_ready(bb_for_body3418_io_Out_6_ready),
    .io_Out_6_valid(bb_for_body3418_io_Out_6_valid),
    .io_Out_6_bits_taskID(bb_for_body3418_io_Out_6_bits_taskID),
    .io_Out_6_bits_control(bb_for_body3418_io_Out_6_bits_control),
    .io_Out_7_ready(bb_for_body3418_io_Out_7_ready),
    .io_Out_7_valid(bb_for_body3418_io_Out_7_valid),
    .io_Out_7_bits_taskID(bb_for_body3418_io_Out_7_bits_taskID),
    .io_Out_7_bits_control(bb_for_body3418_io_Out_7_bits_control),
    .io_Out_8_ready(bb_for_body3418_io_Out_8_ready),
    .io_Out_8_valid(bb_for_body3418_io_Out_8_valid),
    .io_Out_8_bits_taskID(bb_for_body3418_io_Out_8_bits_taskID),
    .io_Out_9_ready(bb_for_body3418_io_Out_9_ready),
    .io_Out_9_valid(bb_for_body3418_io_Out_9_valid),
    .io_Out_9_bits_taskID(bb_for_body3418_io_Out_9_bits_taskID),
    .io_Out_9_bits_control(bb_for_body3418_io_Out_9_bits_control),
    .io_Out_10_ready(bb_for_body3418_io_Out_10_ready),
    .io_Out_10_valid(bb_for_body3418_io_Out_10_valid),
    .io_Out_10_bits_taskID(bb_for_body3418_io_Out_10_bits_taskID),
    .io_Out_10_bits_control(bb_for_body3418_io_Out_10_bits_control),
    .io_Out_11_ready(bb_for_body3418_io_Out_11_ready),
    .io_Out_11_valid(bb_for_body3418_io_Out_11_valid),
    .io_Out_11_bits_taskID(bb_for_body3418_io_Out_11_bits_taskID),
    .io_Out_11_bits_control(bb_for_body3418_io_Out_11_bits_control),
    .io_Out_12_ready(bb_for_body3418_io_Out_12_ready),
    .io_Out_12_valid(bb_for_body3418_io_Out_12_valid),
    .io_Out_12_bits_taskID(bb_for_body3418_io_Out_12_bits_taskID),
    .io_Out_12_bits_control(bb_for_body3418_io_Out_12_bits_control),
    .io_predicateIn_0_ready(bb_for_body3418_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body3418_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body3418_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body3418_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body3418_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body3418_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body3418_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body3418_io_predicateIn_1_bits_control)
  );
  ComputeNode binaryOp_add0 ( // @[extracted_function_reduction.scala 125:29]
    .clock(binaryOp_add0_clock),
    .reset(binaryOp_add0_reset),
    .io_enable_ready(binaryOp_add0_io_enable_ready),
    .io_enable_valid(binaryOp_add0_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add0_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add0_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add0_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add0_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add0_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add0_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add0_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add0_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add0_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add0_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add0_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add0_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add0_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add0_io_RightIO_bits_data)
  );
  ComputeNode_1 icmp_cmp1421 ( // @[extracted_function_reduction.scala 128:28]
    .clock(icmp_cmp1421_clock),
    .reset(icmp_cmp1421_reset),
    .io_enable_ready(icmp_cmp1421_io_enable_ready),
    .io_enable_valid(icmp_cmp1421_io_enable_valid),
    .io_enable_bits_taskID(icmp_cmp1421_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_cmp1421_io_enable_bits_control),
    .io_Out_0_ready(icmp_cmp1421_io_Out_0_ready),
    .io_Out_0_valid(icmp_cmp1421_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_cmp1421_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_cmp1421_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_cmp1421_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_cmp1421_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_cmp1421_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_cmp1421_io_RightIO_ready),
    .io_RightIO_valid(icmp_cmp1421_io_RightIO_valid),
    .io_RightIO_bits_data(icmp_cmp1421_io_RightIO_bits_data)
  );
  CBranchNodeVariable br_2 ( // @[extracted_function_reduction.scala 131:20]
    .clock(br_2_clock),
    .reset(br_2_reset),
    .io_enable_ready(br_2_io_enable_ready),
    .io_enable_valid(br_2_io_enable_valid),
    .io_enable_bits_taskID(br_2_io_enable_bits_taskID),
    .io_enable_bits_control(br_2_io_enable_bits_control),
    .io_CmpIO_ready(br_2_io_CmpIO_ready),
    .io_CmpIO_valid(br_2_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_2_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_2_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_2_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_2_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_2_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_2_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_2_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_2_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_2_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_2_io_FalseOutput_0_bits_control)
  );
  ComputeNode_2 binaryOp_add43 ( // @[extracted_function_reduction.scala 134:30]
    .clock(binaryOp_add43_clock),
    .reset(binaryOp_add43_reset),
    .io_enable_ready(binaryOp_add43_io_enable_ready),
    .io_enable_valid(binaryOp_add43_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add43_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add43_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add43_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add43_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add43_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add43_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add43_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add43_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add43_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add43_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add43_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add43_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add43_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add43_io_RightIO_bits_data)
  );
  ComputeNode_3 icmp_cmp51394 ( // @[extracted_function_reduction.scala 137:29]
    .clock(icmp_cmp51394_clock),
    .reset(icmp_cmp51394_reset),
    .io_enable_ready(icmp_cmp51394_io_enable_ready),
    .io_enable_valid(icmp_cmp51394_io_enable_valid),
    .io_enable_bits_taskID(icmp_cmp51394_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_cmp51394_io_enable_bits_control),
    .io_Out_0_ready(icmp_cmp51394_io_Out_0_ready),
    .io_Out_0_valid(icmp_cmp51394_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_cmp51394_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_cmp51394_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_cmp51394_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_cmp51394_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_cmp51394_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_cmp51394_io_RightIO_ready),
    .io_RightIO_valid(icmp_cmp51394_io_RightIO_valid),
    .io_RightIO_bits_data(icmp_cmp51394_io_RightIO_bits_data)
  );
  ComputeNode_4 binaryOp_add125 ( // @[extracted_function_reduction.scala 140:31]
    .clock(binaryOp_add125_clock),
    .reset(binaryOp_add125_reset),
    .io_enable_ready(binaryOp_add125_io_enable_ready),
    .io_enable_valid(binaryOp_add125_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add125_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add125_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add125_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add125_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add125_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add125_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add125_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add125_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add125_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add125_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add125_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add125_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add125_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add125_io_RightIO_bits_data)
  );
  ComputeNode_5 icmp_cmp131376 ( // @[extracted_function_reduction.scala 143:30]
    .clock(icmp_cmp131376_clock),
    .reset(icmp_cmp131376_reset),
    .io_enable_ready(icmp_cmp131376_io_enable_ready),
    .io_enable_valid(icmp_cmp131376_io_enable_valid),
    .io_enable_bits_taskID(icmp_cmp131376_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_cmp131376_io_enable_bits_control),
    .io_Out_0_ready(icmp_cmp131376_io_Out_0_ready),
    .io_Out_0_valid(icmp_cmp131376_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_cmp131376_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_cmp131376_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_cmp131376_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_cmp131376_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_cmp131376_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_cmp131376_io_RightIO_ready),
    .io_RightIO_valid(icmp_cmp131376_io_RightIO_valid),
    .io_RightIO_bits_data(icmp_cmp131376_io_RightIO_bits_data)
  );
  UBranchNode br_7 ( // @[extracted_function_reduction.scala 146:20]
    .clock(br_7_clock),
    .reset(br_7_reset),
    .io_enable_ready(br_7_io_enable_ready),
    .io_enable_valid(br_7_io_enable_valid),
    .io_enable_bits_taskID(br_7_io_enable_bits_taskID),
    .io_enable_bits_control(br_7_io_enable_bits_control),
    .io_Out_0_ready(br_7_io_Out_0_ready),
    .io_Out_0_valid(br_7_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_7_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_7_io_Out_0_bits_control)
  );
  UBranchNode_1 br_8 ( // @[extracted_function_reduction.scala 149:20]
    .clock(br_8_clock),
    .reset(br_8_reset),
    .io_enable_ready(br_8_io_enable_ready),
    .io_enable_valid(br_8_io_enable_valid),
    .io_enable_bits_taskID(br_8_io_enable_bits_taskID),
    .io_enable_bits_control(br_8_io_enable_bits_control),
    .io_Out_0_ready(br_8_io_Out_0_ready),
    .io_Out_0_valid(br_8_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_8_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_8_io_Out_0_bits_control)
  );
  RetNode2 ret_9 ( // @[extracted_function_reduction.scala 152:21]
    .clock(ret_9_clock),
    .reset(ret_9_reset),
    .io_In_enable_ready(ret_9_io_In_enable_ready),
    .io_In_enable_valid(ret_9_io_In_enable_valid),
    .io_In_enable_bits_taskID(ret_9_io_In_enable_bits_taskID),
    .io_In_enable_bits_control(ret_9_io_In_enable_bits_control),
    .io_Out_ready(ret_9_io_Out_ready),
    .io_Out_valid(ret_9_io_Out_valid),
    .io_Out_bits_enable_taskID(ret_9_io_Out_bits_enable_taskID),
    .io_Out_bits_enable_control(ret_9_io_Out_bits_enable_control)
  );
  PhiFastNode phi_pw_conv_reduction_s1_k_014310 ( // @[extracted_function_reduction.scala 155:49]
    .clock(phi_pw_conv_reduction_s1_k_014310_clock),
    .reset(phi_pw_conv_reduction_s1_k_014310_reset),
    .io_enable_ready(phi_pw_conv_reduction_s1_k_014310_io_enable_ready),
    .io_enable_valid(phi_pw_conv_reduction_s1_k_014310_io_enable_valid),
    .io_enable_bits_control(phi_pw_conv_reduction_s1_k_014310_io_enable_bits_control),
    .io_InData_0_ready(phi_pw_conv_reduction_s1_k_014310_io_InData_0_ready),
    .io_InData_0_valid(phi_pw_conv_reduction_s1_k_014310_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_pw_conv_reduction_s1_k_014310_io_InData_0_bits_taskID),
    .io_InData_0_bits_data(phi_pw_conv_reduction_s1_k_014310_io_InData_0_bits_data),
    .io_InData_1_ready(phi_pw_conv_reduction_s1_k_014310_io_InData_1_ready),
    .io_InData_1_valid(phi_pw_conv_reduction_s1_k_014310_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_pw_conv_reduction_s1_k_014310_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_pw_conv_reduction_s1_k_014310_io_InData_1_bits_data),
    .io_Mask_ready(phi_pw_conv_reduction_s1_k_014310_io_Mask_ready),
    .io_Mask_valid(phi_pw_conv_reduction_s1_k_014310_io_Mask_valid),
    .io_Mask_bits(phi_pw_conv_reduction_s1_k_014310_io_Mask_bits),
    .io_Out_0_ready(phi_pw_conv_reduction_s1_k_014310_io_Out_0_ready),
    .io_Out_0_valid(phi_pw_conv_reduction_s1_k_014310_io_Out_0_valid),
    .io_Out_0_bits_data(phi_pw_conv_reduction_s1_k_014310_io_Out_0_bits_data),
    .io_Out_1_ready(phi_pw_conv_reduction_s1_k_014310_io_Out_1_ready),
    .io_Out_1_valid(phi_pw_conv_reduction_s1_k_014310_io_Out_1_valid),
    .io_Out_1_bits_data(phi_pw_conv_reduction_s1_k_014310_io_Out_1_bits_data)
  );
  ComputeNode_6 binaryOp_sub11 ( // @[extracted_function_reduction.scala 158:30]
    .clock(binaryOp_sub11_clock),
    .reset(binaryOp_sub11_reset),
    .io_enable_ready(binaryOp_sub11_io_enable_ready),
    .io_enable_valid(binaryOp_sub11_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_sub11_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_sub11_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_sub11_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_sub11_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_sub11_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_sub11_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_sub11_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_sub11_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_sub11_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_sub11_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_sub11_io_RightIO_bits_data)
  );
  ComputeNode_7 binaryOp_mul112 ( // @[extracted_function_reduction.scala 161:31]
    .clock(binaryOp_mul112_clock),
    .reset(binaryOp_mul112_reset),
    .io_enable_ready(binaryOp_mul112_io_enable_ready),
    .io_enable_valid(binaryOp_mul112_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul112_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul112_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul112_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul112_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul112_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul112_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul112_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul112_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul112_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul112_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul112_io_RightIO_bits_data)
  );
  CBranchNodeVariable_1 br_13 ( // @[extracted_function_reduction.scala 164:21]
    .clock(br_13_clock),
    .reset(br_13_reset),
    .io_enable_ready(br_13_io_enable_ready),
    .io_enable_valid(br_13_io_enable_valid),
    .io_enable_bits_taskID(br_13_io_enable_bits_taskID),
    .io_enable_bits_control(br_13_io_enable_bits_control),
    .io_CmpIO_ready(br_13_io_CmpIO_ready),
    .io_CmpIO_valid(br_13_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_13_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_13_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_13_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_13_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_13_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_13_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_13_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_13_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_13_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_13_io_FalseOutput_0_bits_control)
  );
  UBranchNode_2 br_14 ( // @[extracted_function_reduction.scala 167:21]
    .clock(br_14_clock),
    .reset(br_14_reset),
    .io_enable_ready(br_14_io_enable_ready),
    .io_enable_valid(br_14_io_enable_valid),
    .io_enable_bits_taskID(br_14_io_enable_bits_taskID),
    .io_enable_bits_control(br_14_io_enable_bits_control),
    .io_Out_0_ready(br_14_io_Out_0_ready),
    .io_Out_0_valid(br_14_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_14_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_14_io_Out_0_bits_control)
  );
  UBranchNode_3 br_15 ( // @[extracted_function_reduction.scala 170:21]
    .clock(br_15_clock),
    .reset(br_15_reset),
    .io_enable_ready(br_15_io_enable_ready),
    .io_enable_valid(br_15_io_enable_valid),
    .io_enable_bits_taskID(br_15_io_enable_bits_taskID),
    .io_enable_bits_control(br_15_io_enable_bits_control),
    .io_Out_0_ready(br_15_io_Out_0_ready),
    .io_Out_0_valid(br_15_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_15_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_15_io_Out_0_bits_control)
  );
  ComputeNode_8 binaryOp_inc6416 ( // @[extracted_function_reduction.scala 173:32]
    .clock(binaryOp_inc6416_clock),
    .reset(binaryOp_inc6416_reset),
    .io_enable_ready(binaryOp_inc6416_io_enable_ready),
    .io_enable_valid(binaryOp_inc6416_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_inc6416_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_inc6416_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_inc6416_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_inc6416_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_inc6416_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_inc6416_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_inc6416_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_inc6416_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_inc6416_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_inc6416_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_inc6416_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_inc6416_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_inc6416_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_inc6416_io_RightIO_valid)
  );
  ComputeNode_9 icmp_exitcond14817 ( // @[extracted_function_reduction.scala 176:34]
    .clock(icmp_exitcond14817_clock),
    .reset(icmp_exitcond14817_reset),
    .io_enable_ready(icmp_exitcond14817_io_enable_ready),
    .io_enable_valid(icmp_exitcond14817_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond14817_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond14817_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond14817_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond14817_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond14817_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond14817_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond14817_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond14817_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond14817_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond14817_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond14817_io_RightIO_valid),
    .io_RightIO_bits_data(icmp_exitcond14817_io_RightIO_bits_data)
  );
  CBranchNodeVariable_2 br_18 ( // @[extracted_function_reduction.scala 179:21]
    .clock(br_18_clock),
    .reset(br_18_reset),
    .io_enable_ready(br_18_io_enable_ready),
    .io_enable_valid(br_18_io_enable_valid),
    .io_enable_bits_taskID(br_18_io_enable_bits_taskID),
    .io_enable_bits_control(br_18_io_enable_bits_control),
    .io_CmpIO_ready(br_18_io_CmpIO_ready),
    .io_CmpIO_valid(br_18_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_18_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_18_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_18_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_18_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_18_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_18_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_18_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_18_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_18_io_FalseOutput_0_bits_control)
  );
  PhiFastNode_1 phi_pw_conv_reduction_s1_y_014019 ( // @[extracted_function_reduction.scala 182:49]
    .clock(phi_pw_conv_reduction_s1_y_014019_clock),
    .reset(phi_pw_conv_reduction_s1_y_014019_reset),
    .io_enable_ready(phi_pw_conv_reduction_s1_y_014019_io_enable_ready),
    .io_enable_valid(phi_pw_conv_reduction_s1_y_014019_io_enable_valid),
    .io_enable_bits_control(phi_pw_conv_reduction_s1_y_014019_io_enable_bits_control),
    .io_InData_0_ready(phi_pw_conv_reduction_s1_y_014019_io_InData_0_ready),
    .io_InData_0_valid(phi_pw_conv_reduction_s1_y_014019_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_pw_conv_reduction_s1_y_014019_io_InData_0_bits_taskID),
    .io_InData_0_bits_data(phi_pw_conv_reduction_s1_y_014019_io_InData_0_bits_data),
    .io_InData_1_ready(phi_pw_conv_reduction_s1_y_014019_io_InData_1_ready),
    .io_InData_1_valid(phi_pw_conv_reduction_s1_y_014019_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_pw_conv_reduction_s1_y_014019_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_pw_conv_reduction_s1_y_014019_io_InData_1_bits_data),
    .io_Mask_ready(phi_pw_conv_reduction_s1_y_014019_io_Mask_ready),
    .io_Mask_valid(phi_pw_conv_reduction_s1_y_014019_io_Mask_valid),
    .io_Mask_bits(phi_pw_conv_reduction_s1_y_014019_io_Mask_bits),
    .io_Out_0_ready(phi_pw_conv_reduction_s1_y_014019_io_Out_0_ready),
    .io_Out_0_valid(phi_pw_conv_reduction_s1_y_014019_io_Out_0_valid),
    .io_Out_0_bits_data(phi_pw_conv_reduction_s1_y_014019_io_Out_0_bits_data),
    .io_Out_1_ready(phi_pw_conv_reduction_s1_y_014019_io_Out_1_ready),
    .io_Out_1_valid(phi_pw_conv_reduction_s1_y_014019_io_Out_1_valid),
    .io_Out_1_bits_data(phi_pw_conv_reduction_s1_y_014019_io_Out_1_bits_data),
    .io_Out_2_ready(phi_pw_conv_reduction_s1_y_014019_io_Out_2_ready),
    .io_Out_2_valid(phi_pw_conv_reduction_s1_y_014019_io_Out_2_valid),
    .io_Out_2_bits_data(phi_pw_conv_reduction_s1_y_014019_io_Out_2_bits_data)
  );
  CBranchNodeVariable_3 br_20 ( // @[extracted_function_reduction.scala 185:21]
    .clock(br_20_clock),
    .reset(br_20_reset),
    .io_enable_ready(br_20_io_enable_ready),
    .io_enable_valid(br_20_io_enable_valid),
    .io_enable_bits_taskID(br_20_io_enable_bits_taskID),
    .io_enable_bits_control(br_20_io_enable_bits_control),
    .io_CmpIO_ready(br_20_io_CmpIO_ready),
    .io_CmpIO_valid(br_20_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_20_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_20_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_20_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_20_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_taskID(br_20_io_TrueOutput_0_bits_taskID),
    .io_TrueOutput_0_bits_control(br_20_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_20_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_20_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_20_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_20_io_FalseOutput_0_bits_control)
  );
  ComputeNode_10 binaryOp_sub821 ( // @[extracted_function_reduction.scala 188:31]
    .clock(binaryOp_sub821_clock),
    .reset(binaryOp_sub821_reset),
    .io_enable_ready(binaryOp_sub821_io_enable_ready),
    .io_enable_valid(binaryOp_sub821_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_sub821_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_sub821_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_sub821_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_sub821_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_sub821_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_sub821_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_sub821_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_sub821_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_sub821_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_sub821_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_sub821_io_RightIO_bits_data)
  );
  ComputeNode_11 binaryOp_reass_add22 ( // @[extracted_function_reduction.scala 191:36]
    .clock(binaryOp_reass_add22_clock),
    .reset(binaryOp_reass_add22_reset),
    .io_enable_ready(binaryOp_reass_add22_io_enable_ready),
    .io_enable_valid(binaryOp_reass_add22_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_reass_add22_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_reass_add22_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_reass_add22_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_reass_add22_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_reass_add22_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_reass_add22_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_reass_add22_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_reass_add22_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_reass_add22_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_reass_add22_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_reass_add22_io_RightIO_bits_data)
  );
  ComputeNode_12 binaryOp_reass_mul23 ( // @[extracted_function_reduction.scala 194:36]
    .clock(binaryOp_reass_mul23_clock),
    .reset(binaryOp_reass_mul23_reset),
    .io_enable_ready(binaryOp_reass_mul23_io_enable_ready),
    .io_enable_valid(binaryOp_reass_mul23_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_reass_mul23_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_reass_mul23_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_reass_mul23_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_reass_mul23_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_reass_mul23_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_reass_mul23_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_reass_mul23_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_reass_mul23_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_reass_mul23_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_reass_mul23_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_reass_mul23_io_RightIO_bits_data)
  );
  UBranchNode_4 br_24 ( // @[extracted_function_reduction.scala 197:21]
    .clock(br_24_clock),
    .reset(br_24_reset),
    .io_enable_ready(br_24_io_enable_ready),
    .io_enable_valid(br_24_io_enable_valid),
    .io_enable_bits_taskID(br_24_io_enable_bits_taskID),
    .io_enable_bits_control(br_24_io_enable_bits_control),
    .io_Out_0_ready(br_24_io_Out_0_ready),
    .io_Out_0_valid(br_24_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_24_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_24_io_Out_0_bits_control)
  );
  UBranchNode_5 br_25 ( // @[extracted_function_reduction.scala 200:21]
    .clock(br_25_clock),
    .reset(br_25_reset),
    .io_enable_ready(br_25_io_enable_ready),
    .io_enable_valid(br_25_io_enable_valid),
    .io_enable_bits_taskID(br_25_io_enable_bits_taskID),
    .io_enable_bits_control(br_25_io_enable_bits_control),
    .io_Out_0_ready(br_25_io_Out_0_ready),
    .io_Out_0_valid(br_25_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_25_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_25_io_Out_0_bits_control)
  );
  ComputeNode_13 binaryOp_inc6126 ( // @[extracted_function_reduction.scala 203:32]
    .clock(binaryOp_inc6126_clock),
    .reset(binaryOp_inc6126_reset),
    .io_enable_ready(binaryOp_inc6126_io_enable_ready),
    .io_enable_valid(binaryOp_inc6126_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_inc6126_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_inc6126_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_inc6126_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_inc6126_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_inc6126_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_inc6126_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_inc6126_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_inc6126_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_inc6126_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_inc6126_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_inc6126_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_inc6126_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_inc6126_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_inc6126_io_RightIO_valid)
  );
  ComputeNode_14 icmp_exitcond14727 ( // @[extracted_function_reduction.scala 206:34]
    .clock(icmp_exitcond14727_clock),
    .reset(icmp_exitcond14727_reset),
    .io_enable_ready(icmp_exitcond14727_io_enable_ready),
    .io_enable_valid(icmp_exitcond14727_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond14727_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond14727_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond14727_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond14727_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond14727_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond14727_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond14727_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond14727_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond14727_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond14727_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond14727_io_RightIO_valid),
    .io_RightIO_bits_data(icmp_exitcond14727_io_RightIO_bits_data)
  );
  CBranchNodeVariable_4 br_28 ( // @[extracted_function_reduction.scala 209:21]
    .clock(br_28_clock),
    .reset(br_28_reset),
    .io_enable_ready(br_28_io_enable_ready),
    .io_enable_valid(br_28_io_enable_valid),
    .io_enable_bits_taskID(br_28_io_enable_bits_taskID),
    .io_enable_bits_control(br_28_io_enable_bits_control),
    .io_CmpIO_ready(br_28_io_CmpIO_ready),
    .io_CmpIO_valid(br_28_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_28_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_28_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_28_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_28_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_28_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_28_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_28_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_28_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_28_io_FalseOutput_0_bits_control)
  );
  PhiFastNode_2 phi_pw_conv_reduction_s1_x_013829 ( // @[extracted_function_reduction.scala 212:49]
    .clock(phi_pw_conv_reduction_s1_x_013829_clock),
    .reset(phi_pw_conv_reduction_s1_x_013829_reset),
    .io_enable_ready(phi_pw_conv_reduction_s1_x_013829_io_enable_ready),
    .io_enable_valid(phi_pw_conv_reduction_s1_x_013829_io_enable_valid),
    .io_enable_bits_control(phi_pw_conv_reduction_s1_x_013829_io_enable_bits_control),
    .io_InData_0_ready(phi_pw_conv_reduction_s1_x_013829_io_InData_0_ready),
    .io_InData_0_valid(phi_pw_conv_reduction_s1_x_013829_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_pw_conv_reduction_s1_x_013829_io_InData_0_bits_taskID),
    .io_InData_0_bits_data(phi_pw_conv_reduction_s1_x_013829_io_InData_0_bits_data),
    .io_InData_1_ready(phi_pw_conv_reduction_s1_x_013829_io_InData_1_ready),
    .io_InData_1_valid(phi_pw_conv_reduction_s1_x_013829_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_pw_conv_reduction_s1_x_013829_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_pw_conv_reduction_s1_x_013829_io_InData_1_bits_data),
    .io_Mask_ready(phi_pw_conv_reduction_s1_x_013829_io_Mask_ready),
    .io_Mask_valid(phi_pw_conv_reduction_s1_x_013829_io_Mask_valid),
    .io_Mask_bits(phi_pw_conv_reduction_s1_x_013829_io_Mask_bits),
    .io_Out_0_ready(phi_pw_conv_reduction_s1_x_013829_io_Out_0_ready),
    .io_Out_0_valid(phi_pw_conv_reduction_s1_x_013829_io_Out_0_valid),
    .io_Out_0_bits_data(phi_pw_conv_reduction_s1_x_013829_io_Out_0_bits_data),
    .io_Out_1_ready(phi_pw_conv_reduction_s1_x_013829_io_Out_1_ready),
    .io_Out_1_valid(phi_pw_conv_reduction_s1_x_013829_io_Out_1_valid),
    .io_Out_1_bits_data(phi_pw_conv_reduction_s1_x_013829_io_Out_1_bits_data),
    .io_Out_2_ready(phi_pw_conv_reduction_s1_x_013829_io_Out_2_ready),
    .io_Out_2_valid(phi_pw_conv_reduction_s1_x_013829_io_Out_2_valid),
    .io_Out_2_bits_data(phi_pw_conv_reduction_s1_x_013829_io_Out_2_bits_data)
  );
  ComputeNode_15 binaryOp_sub1630 ( // @[extracted_function_reduction.scala 215:32]
    .clock(binaryOp_sub1630_clock),
    .reset(binaryOp_sub1630_reset),
    .io_enable_ready(binaryOp_sub1630_io_enable_ready),
    .io_enable_valid(binaryOp_sub1630_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_sub1630_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_sub1630_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_sub1630_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_sub1630_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_sub1630_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_sub1630_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_sub1630_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_sub1630_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_sub1630_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_sub1630_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_sub1630_io_RightIO_bits_data)
  );
  ComputeNode_16 binaryOp_add1031 ( // @[extracted_function_reduction.scala 218:32]
    .clock(binaryOp_add1031_clock),
    .reset(binaryOp_add1031_reset),
    .io_enable_ready(binaryOp_add1031_io_enable_ready),
    .io_enable_valid(binaryOp_add1031_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add1031_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add1031_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add1031_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add1031_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add1031_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add1031_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add1031_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add1031_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add1031_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add1031_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add1031_io_RightIO_bits_data)
  );
  ComputeNode_17 binaryOp_add1732 ( // @[extracted_function_reduction.scala 221:32]
    .clock(binaryOp_add1732_clock),
    .reset(binaryOp_add1732_reset),
    .io_enable_ready(binaryOp_add1732_io_enable_ready),
    .io_enable_valid(binaryOp_add1732_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add1732_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add1732_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add1732_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add1732_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add1732_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add1732_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add1732_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add1732_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add1732_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add1732_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add1732_io_RightIO_bits_data)
  );
  GepNode Gep_arrayidx5033 ( // @[extracted_function_reduction.scala 224:32]
    .clock(Gep_arrayidx5033_clock),
    .reset(Gep_arrayidx5033_reset),
    .io_enable_ready(Gep_arrayidx5033_io_enable_ready),
    .io_enable_valid(Gep_arrayidx5033_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx5033_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx5033_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx5033_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx5033_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx5033_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx5033_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx5033_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx5033_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx5033_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx5033_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx5033_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx5033_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx5033_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx5033_io_idx_0_bits_data)
  );
  UBranchNode_6 br_34 ( // @[extracted_function_reduction.scala 227:21]
    .clock(br_34_clock),
    .reset(br_34_reset),
    .io_enable_ready(br_34_io_enable_ready),
    .io_enable_valid(br_34_io_enable_valid),
    .io_enable_bits_taskID(br_34_io_enable_bits_taskID),
    .io_enable_bits_control(br_34_io_enable_bits_control),
    .io_Out_0_ready(br_34_io_Out_0_ready),
    .io_Out_0_valid(br_34_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_34_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_34_io_Out_0_bits_control)
  );
  ComputeNode_18 binaryOp_inc5835 ( // @[extracted_function_reduction.scala 230:32]
    .clock(binaryOp_inc5835_clock),
    .reset(binaryOp_inc5835_reset),
    .io_enable_ready(binaryOp_inc5835_io_enable_ready),
    .io_enable_valid(binaryOp_inc5835_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_inc5835_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_inc5835_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_inc5835_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_inc5835_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_inc5835_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_inc5835_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_inc5835_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_inc5835_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_inc5835_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_inc5835_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_inc5835_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_inc5835_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_inc5835_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_inc5835_io_RightIO_valid)
  );
  ComputeNode_19 icmp_exitcond14636 ( // @[extracted_function_reduction.scala 233:34]
    .clock(icmp_exitcond14636_clock),
    .reset(icmp_exitcond14636_reset),
    .io_enable_ready(icmp_exitcond14636_io_enable_ready),
    .io_enable_valid(icmp_exitcond14636_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond14636_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond14636_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond14636_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond14636_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond14636_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond14636_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond14636_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond14636_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond14636_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond14636_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond14636_io_RightIO_valid),
    .io_RightIO_bits_data(icmp_exitcond14636_io_RightIO_bits_data)
  );
  CBranchNodeVariable_5 br_37 ( // @[extracted_function_reduction.scala 236:21]
    .clock(br_37_clock),
    .reset(br_37_reset),
    .io_enable_ready(br_37_io_enable_ready),
    .io_enable_valid(br_37_io_enable_valid),
    .io_enable_bits_taskID(br_37_io_enable_bits_taskID),
    .io_enable_bits_control(br_37_io_enable_bits_control),
    .io_CmpIO_ready(br_37_io_CmpIO_ready),
    .io_CmpIO_valid(br_37_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_37_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_37_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_37_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_37_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_37_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_37_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_37_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_37_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_37_io_FalseOutput_0_bits_control)
  );
  PhiFastNode_3 phi_pw_conv_reduction_s1_r_pw__x_013638 ( // @[extracted_function_reduction.scala 239:55]
    .clock(phi_pw_conv_reduction_s1_r_pw__x_013638_clock),
    .reset(phi_pw_conv_reduction_s1_r_pw__x_013638_reset),
    .io_enable_ready(phi_pw_conv_reduction_s1_r_pw__x_013638_io_enable_ready),
    .io_enable_valid(phi_pw_conv_reduction_s1_r_pw__x_013638_io_enable_valid),
    .io_enable_bits_control(phi_pw_conv_reduction_s1_r_pw__x_013638_io_enable_bits_control),
    .io_InData_0_ready(phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_0_ready),
    .io_InData_0_valid(phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_ready),
    .io_InData_1_valid(phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_bits_data),
    .io_Mask_ready(phi_pw_conv_reduction_s1_r_pw__x_013638_io_Mask_ready),
    .io_Mask_valid(phi_pw_conv_reduction_s1_r_pw__x_013638_io_Mask_valid),
    .io_Mask_bits(phi_pw_conv_reduction_s1_r_pw__x_013638_io_Mask_bits),
    .io_Out_0_ready(phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_0_ready),
    .io_Out_0_valid(phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_0_valid),
    .io_Out_0_bits_data(phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_0_bits_data),
    .io_Out_1_ready(phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_1_ready),
    .io_Out_1_valid(phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_1_valid),
    .io_Out_1_bits_data(phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_1_bits_data)
  );
  ComputeNode_20 binaryOp_mul2239 ( // @[extracted_function_reduction.scala 242:32]
    .clock(binaryOp_mul2239_clock),
    .reset(binaryOp_mul2239_reset),
    .io_enable_ready(binaryOp_mul2239_io_enable_ready),
    .io_enable_valid(binaryOp_mul2239_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul2239_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul2239_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul2239_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul2239_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul2239_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul2239_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul2239_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul2239_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul2239_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul2239_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul2239_io_RightIO_bits_data)
  );
  ComputeNode_21 binaryOp_add2340 ( // @[extracted_function_reduction.scala 245:32]
    .clock(binaryOp_add2340_clock),
    .reset(binaryOp_add2340_reset),
    .io_enable_ready(binaryOp_add2340_io_enable_ready),
    .io_enable_valid(binaryOp_add2340_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add2340_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add2340_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add2340_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add2340_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add2340_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add2340_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add2340_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add2340_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add2340_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add2340_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add2340_io_RightIO_bits_data)
  );
  UBranchNode_7 br_41 ( // @[extracted_function_reduction.scala 248:21]
    .clock(br_41_clock),
    .reset(br_41_reset),
    .io_enable_ready(br_41_io_enable_ready),
    .io_enable_valid(br_41_io_enable_valid),
    .io_enable_bits_taskID(br_41_io_enable_bits_taskID),
    .io_enable_bits_control(br_41_io_enable_bits_control),
    .io_Out_0_ready(br_41_io_Out_0_ready),
    .io_Out_0_valid(br_41_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_41_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_41_io_Out_0_bits_control)
  );
  PhiFastNode_4 phiadd38_lcssa_lcssa42 ( // @[extracted_function_reduction.scala 251:38]
    .clock(phiadd38_lcssa_lcssa42_clock),
    .reset(phiadd38_lcssa_lcssa42_reset),
    .io_enable_ready(phiadd38_lcssa_lcssa42_io_enable_ready),
    .io_enable_valid(phiadd38_lcssa_lcssa42_io_enable_valid),
    .io_enable_bits_control(phiadd38_lcssa_lcssa42_io_enable_bits_control),
    .io_InData_0_ready(phiadd38_lcssa_lcssa42_io_InData_0_ready),
    .io_InData_0_valid(phiadd38_lcssa_lcssa42_io_InData_0_valid),
    .io_InData_0_bits_taskID(phiadd38_lcssa_lcssa42_io_InData_0_bits_taskID),
    .io_InData_0_bits_data(phiadd38_lcssa_lcssa42_io_InData_0_bits_data),
    .io_Out_0_ready(phiadd38_lcssa_lcssa42_io_Out_0_ready),
    .io_Out_0_valid(phiadd38_lcssa_lcssa42_io_Out_0_valid),
    .io_Out_0_bits_data(phiadd38_lcssa_lcssa42_io_Out_0_bits_data)
  );
  ComputeNode_22 binaryOp_mul4443 ( // @[extracted_function_reduction.scala 254:32]
    .clock(binaryOp_mul4443_clock),
    .reset(binaryOp_mul4443_reset),
    .io_enable_ready(binaryOp_mul4443_io_enable_ready),
    .io_enable_valid(binaryOp_mul4443_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul4443_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul4443_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul4443_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul4443_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul4443_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul4443_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul4443_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul4443_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul4443_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul4443_io_RightIO_valid)
  );
  SextNode sextconv4744 ( // @[extracted_function_reduction.scala 257:28]
    .clock(sextconv4744_clock),
    .reset(sextconv4744_reset),
    .io_Input_ready(sextconv4744_io_Input_ready),
    .io_Input_valid(sextconv4744_io_Input_valid),
    .io_Input_bits_data(sextconv4744_io_Input_bits_data),
    .io_enable_ready(sextconv4744_io_enable_ready),
    .io_enable_valid(sextconv4744_io_enable_valid),
    .io_enable_bits_taskID(sextconv4744_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv4744_io_Out_0_ready),
    .io_Out_0_valid(sextconv4744_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv4744_io_Out_0_bits_data)
  );
  UnTypLoad ld_45 ( // @[extracted_function_reduction.scala 260:21]
    .clock(ld_45_clock),
    .reset(ld_45_reset),
    .io_enable_ready(ld_45_io_enable_ready),
    .io_enable_valid(ld_45_io_enable_valid),
    .io_enable_bits_taskID(ld_45_io_enable_bits_taskID),
    .io_enable_bits_control(ld_45_io_enable_bits_control),
    .io_Out_0_ready(ld_45_io_Out_0_ready),
    .io_Out_0_valid(ld_45_io_Out_0_valid),
    .io_Out_0_bits_data(ld_45_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_45_io_GepAddr_ready),
    .io_GepAddr_valid(ld_45_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_45_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_45_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_45_io_GepAddr_bits_data),
    .io_memReq_ready(ld_45_io_memReq_ready),
    .io_memReq_valid(ld_45_io_memReq_valid),
    .io_memReq_bits_address(ld_45_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_45_io_memReq_bits_taskID),
    .io_memResp_valid(ld_45_io_memResp_valid),
    .io_memResp_data(ld_45_io_memResp_data)
  );
  ComputeNode_23 binaryOp_add5246 ( // @[extracted_function_reduction.scala 263:32]
    .clock(binaryOp_add5246_clock),
    .reset(binaryOp_add5246_reset),
    .io_enable_ready(binaryOp_add5246_io_enable_ready),
    .io_enable_valid(binaryOp_add5246_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add5246_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add5246_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add5246_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add5246_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add5246_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add5246_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add5246_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add5246_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add5246_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add5246_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add5246_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add5246_io_RightIO_bits_data)
  );
  UnTypStore st_47 ( // @[extracted_function_reduction.scala 266:21]
    .clock(st_47_clock),
    .reset(st_47_reset),
    .io_enable_ready(st_47_io_enable_ready),
    .io_enable_valid(st_47_io_enable_valid),
    .io_enable_bits_taskID(st_47_io_enable_bits_taskID),
    .io_enable_bits_control(st_47_io_enable_bits_control),
    .io_GepAddr_ready(st_47_io_GepAddr_ready),
    .io_GepAddr_valid(st_47_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_47_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_47_io_GepAddr_bits_data),
    .io_inData_ready(st_47_io_inData_ready),
    .io_inData_valid(st_47_io_inData_valid),
    .io_inData_bits_taskID(st_47_io_inData_bits_taskID),
    .io_inData_bits_data(st_47_io_inData_bits_data),
    .io_memReq_ready(st_47_io_memReq_ready),
    .io_memReq_valid(st_47_io_memReq_valid),
    .io_memReq_bits_address(st_47_io_memReq_bits_address),
    .io_memReq_bits_data(st_47_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_47_io_memReq_bits_taskID),
    .io_memResp_valid(st_47_io_memResp_valid)
  );
  ComputeNode_24 binaryOp_inc5548 ( // @[extracted_function_reduction.scala 269:32]
    .clock(binaryOp_inc5548_clock),
    .reset(binaryOp_inc5548_reset),
    .io_enable_ready(binaryOp_inc5548_io_enable_ready),
    .io_enable_valid(binaryOp_inc5548_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_inc5548_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_inc5548_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_inc5548_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_inc5548_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_inc5548_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_inc5548_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_inc5548_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_inc5548_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_inc5548_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_inc5548_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_inc5548_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_inc5548_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_inc5548_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_inc5548_io_RightIO_valid)
  );
  ComputeNode_25 icmp_exitcond14549 ( // @[extracted_function_reduction.scala 272:34]
    .clock(icmp_exitcond14549_clock),
    .reset(icmp_exitcond14549_reset),
    .io_enable_ready(icmp_exitcond14549_io_enable_ready),
    .io_enable_valid(icmp_exitcond14549_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond14549_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond14549_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond14549_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond14549_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond14549_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond14549_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond14549_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond14549_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond14549_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond14549_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond14549_io_RightIO_valid)
  );
  CBranchNodeVariable_6 br_50 ( // @[extracted_function_reduction.scala 275:21]
    .clock(br_50_clock),
    .reset(br_50_reset),
    .io_enable_ready(br_50_io_enable_ready),
    .io_enable_valid(br_50_io_enable_valid),
    .io_enable_bits_taskID(br_50_io_enable_bits_taskID),
    .io_enable_bits_control(br_50_io_enable_bits_control),
    .io_CmpIO_ready(br_50_io_CmpIO_ready),
    .io_CmpIO_valid(br_50_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_50_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_50_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_50_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_50_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_50_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_50_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_50_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_50_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_50_io_FalseOutput_0_bits_control)
  );
  PhiFastNode_5 phi_dw_conv_013551 ( // @[extracted_function_reduction.scala 278:34]
    .clock(phi_dw_conv_013551_clock),
    .reset(phi_dw_conv_013551_reset),
    .io_enable_ready(phi_dw_conv_013551_io_enable_ready),
    .io_enable_valid(phi_dw_conv_013551_io_enable_valid),
    .io_enable_bits_taskID(phi_dw_conv_013551_io_enable_bits_taskID),
    .io_enable_bits_control(phi_dw_conv_013551_io_enable_bits_control),
    .io_InData_0_ready(phi_dw_conv_013551_io_InData_0_ready),
    .io_InData_0_valid(phi_dw_conv_013551_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_dw_conv_013551_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi_dw_conv_013551_io_InData_1_ready),
    .io_InData_1_valid(phi_dw_conv_013551_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_dw_conv_013551_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_dw_conv_013551_io_InData_1_bits_data),
    .io_Mask_ready(phi_dw_conv_013551_io_Mask_ready),
    .io_Mask_valid(phi_dw_conv_013551_io_Mask_valid),
    .io_Mask_bits(phi_dw_conv_013551_io_Mask_bits),
    .io_Out_0_ready(phi_dw_conv_013551_io_Out_0_ready),
    .io_Out_0_valid(phi_dw_conv_013551_io_Out_0_valid),
    .io_Out_0_bits_taskID(phi_dw_conv_013551_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(phi_dw_conv_013551_io_Out_0_bits_data)
  );
  PhiFastNode_6 phi_dw_conv_s1_r_dw__y_013452 ( // @[extracted_function_reduction.scala 281:45]
    .clock(phi_dw_conv_s1_r_dw__y_013452_clock),
    .reset(phi_dw_conv_s1_r_dw__y_013452_reset),
    .io_enable_ready(phi_dw_conv_s1_r_dw__y_013452_io_enable_ready),
    .io_enable_valid(phi_dw_conv_s1_r_dw__y_013452_io_enable_valid),
    .io_enable_bits_control(phi_dw_conv_s1_r_dw__y_013452_io_enable_bits_control),
    .io_InData_0_ready(phi_dw_conv_s1_r_dw__y_013452_io_InData_0_ready),
    .io_InData_0_valid(phi_dw_conv_s1_r_dw__y_013452_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_dw_conv_s1_r_dw__y_013452_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi_dw_conv_s1_r_dw__y_013452_io_InData_1_ready),
    .io_InData_1_valid(phi_dw_conv_s1_r_dw__y_013452_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_dw_conv_s1_r_dw__y_013452_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_dw_conv_s1_r_dw__y_013452_io_InData_1_bits_data),
    .io_Mask_ready(phi_dw_conv_s1_r_dw__y_013452_io_Mask_ready),
    .io_Mask_valid(phi_dw_conv_s1_r_dw__y_013452_io_Mask_valid),
    .io_Mask_bits(phi_dw_conv_s1_r_dw__y_013452_io_Mask_bits),
    .io_Out_0_ready(phi_dw_conv_s1_r_dw__y_013452_io_Out_0_ready),
    .io_Out_0_valid(phi_dw_conv_s1_r_dw__y_013452_io_Out_0_valid),
    .io_Out_0_bits_data(phi_dw_conv_s1_r_dw__y_013452_io_Out_0_bits_data),
    .io_Out_1_ready(phi_dw_conv_s1_r_dw__y_013452_io_Out_1_ready),
    .io_Out_1_valid(phi_dw_conv_s1_r_dw__y_013452_io_Out_1_valid),
    .io_Out_1_bits_data(phi_dw_conv_s1_r_dw__y_013452_io_Out_1_bits_data)
  );
  ComputeNode_26 binaryOp_add2853 ( // @[extracted_function_reduction.scala 284:32]
    .clock(binaryOp_add2853_clock),
    .reset(binaryOp_add2853_reset),
    .io_enable_ready(binaryOp_add2853_io_enable_ready),
    .io_enable_valid(binaryOp_add2853_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add2853_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add2853_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add2853_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add2853_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add2853_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add2853_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add2853_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add2853_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add2853_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add2853_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add2853_io_RightIO_bits_data)
  );
  ComputeNode_27 binaryOp_mul2954 ( // @[extracted_function_reduction.scala 287:32]
    .clock(binaryOp_mul2954_clock),
    .reset(binaryOp_mul2954_reset),
    .io_enable_ready(binaryOp_mul2954_io_enable_ready),
    .io_enable_valid(binaryOp_mul2954_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul2954_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul2954_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul2954_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul2954_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul2954_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul2954_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul2954_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul2954_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul2954_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul2954_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul2954_io_RightIO_bits_data)
  );
  ComputeNode_28 binaryOp_add3055 ( // @[extracted_function_reduction.scala 290:32]
    .clock(binaryOp_add3055_clock),
    .reset(binaryOp_add3055_reset),
    .io_enable_ready(binaryOp_add3055_io_enable_ready),
    .io_enable_valid(binaryOp_add3055_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add3055_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add3055_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add3055_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add3055_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add3055_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add3055_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add3055_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add3055_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add3055_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add3055_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add3055_io_RightIO_bits_data)
  );
  UBranchNode_8 br_56 ( // @[extracted_function_reduction.scala 293:21]
    .clock(br_56_clock),
    .reset(br_56_reset),
    .io_enable_ready(br_56_io_enable_ready),
    .io_enable_valid(br_56_io_enable_valid),
    .io_enable_bits_taskID(br_56_io_enable_bits_taskID),
    .io_enable_bits_control(br_56_io_enable_bits_control),
    .io_Out_0_ready(br_56_io_Out_0_ready),
    .io_Out_0_valid(br_56_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_56_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_56_io_Out_0_bits_control)
  );
  PhiFastNode_7 phiadd38_lcssa57 ( // @[extracted_function_reduction.scala 296:32]
    .clock(phiadd38_lcssa57_clock),
    .reset(phiadd38_lcssa57_reset),
    .io_enable_ready(phiadd38_lcssa57_io_enable_ready),
    .io_enable_valid(phiadd38_lcssa57_io_enable_valid),
    .io_enable_bits_taskID(phiadd38_lcssa57_io_enable_bits_taskID),
    .io_enable_bits_control(phiadd38_lcssa57_io_enable_bits_control),
    .io_InData_0_ready(phiadd38_lcssa57_io_InData_0_ready),
    .io_InData_0_valid(phiadd38_lcssa57_io_InData_0_valid),
    .io_InData_0_bits_taskID(phiadd38_lcssa57_io_InData_0_bits_taskID),
    .io_InData_0_bits_data(phiadd38_lcssa57_io_InData_0_bits_data),
    .io_Out_0_ready(phiadd38_lcssa57_io_Out_0_ready),
    .io_Out_0_valid(phiadd38_lcssa57_io_Out_0_valid),
    .io_Out_0_bits_taskID(phiadd38_lcssa57_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(phiadd38_lcssa57_io_Out_0_bits_data),
    .io_Out_1_ready(phiadd38_lcssa57_io_Out_1_ready),
    .io_Out_1_valid(phiadd38_lcssa57_io_Out_1_valid),
    .io_Out_1_bits_taskID(phiadd38_lcssa57_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(phiadd38_lcssa57_io_Out_1_bits_data)
  );
  ComputeNode_29 binaryOp_inc4158 ( // @[extracted_function_reduction.scala 299:32]
    .clock(binaryOp_inc4158_clock),
    .reset(binaryOp_inc4158_reset),
    .io_enable_ready(binaryOp_inc4158_io_enable_ready),
    .io_enable_valid(binaryOp_inc4158_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_inc4158_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_inc4158_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_inc4158_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_inc4158_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_inc4158_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_inc4158_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_inc4158_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_inc4158_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_inc4158_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_inc4158_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_inc4158_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_inc4158_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_inc4158_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_inc4158_io_RightIO_valid)
  );
  ComputeNode_30 icmp_exitcond14459 ( // @[extracted_function_reduction.scala 302:34]
    .clock(icmp_exitcond14459_clock),
    .reset(icmp_exitcond14459_reset),
    .io_enable_ready(icmp_exitcond14459_io_enable_ready),
    .io_enable_valid(icmp_exitcond14459_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond14459_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond14459_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond14459_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond14459_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond14459_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond14459_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond14459_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond14459_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond14459_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond14459_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond14459_io_RightIO_valid)
  );
  CBranchNodeVariable_7 br_60 ( // @[extracted_function_reduction.scala 305:21]
    .clock(br_60_clock),
    .reset(br_60_reset),
    .io_enable_ready(br_60_io_enable_ready),
    .io_enable_valid(br_60_io_enable_valid),
    .io_enable_bits_taskID(br_60_io_enable_bits_taskID),
    .io_enable_bits_control(br_60_io_enable_bits_control),
    .io_CmpIO_ready(br_60_io_CmpIO_ready),
    .io_CmpIO_valid(br_60_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_60_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_60_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_60_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_60_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_60_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_60_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_60_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_60_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_60_io_FalseOutput_0_bits_control)
  );
  PhiFastNode_8 phi_dw_conv_113361 ( // @[extracted_function_reduction.scala 308:34]
    .clock(phi_dw_conv_113361_clock),
    .reset(phi_dw_conv_113361_reset),
    .io_enable_ready(phi_dw_conv_113361_io_enable_ready),
    .io_enable_valid(phi_dw_conv_113361_io_enable_valid),
    .io_enable_bits_control(phi_dw_conv_113361_io_enable_bits_control),
    .io_InData_0_ready(phi_dw_conv_113361_io_InData_0_ready),
    .io_InData_0_valid(phi_dw_conv_113361_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_dw_conv_113361_io_InData_0_bits_taskID),
    .io_InData_0_bits_data(phi_dw_conv_113361_io_InData_0_bits_data),
    .io_InData_1_ready(phi_dw_conv_113361_io_InData_1_ready),
    .io_InData_1_valid(phi_dw_conv_113361_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_dw_conv_113361_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_dw_conv_113361_io_InData_1_bits_data),
    .io_Mask_ready(phi_dw_conv_113361_io_Mask_ready),
    .io_Mask_valid(phi_dw_conv_113361_io_Mask_valid),
    .io_Mask_bits(phi_dw_conv_113361_io_Mask_bits),
    .io_Out_0_ready(phi_dw_conv_113361_io_Out_0_ready),
    .io_Out_0_valid(phi_dw_conv_113361_io_Out_0_valid),
    .io_Out_0_bits_data(phi_dw_conv_113361_io_Out_0_bits_data)
  );
  PhiFastNode_9 phi_dw_conv_s1_r_dw__x_013262 ( // @[extracted_function_reduction.scala 311:45]
    .clock(phi_dw_conv_s1_r_dw__x_013262_clock),
    .reset(phi_dw_conv_s1_r_dw__x_013262_reset),
    .io_enable_ready(phi_dw_conv_s1_r_dw__x_013262_io_enable_ready),
    .io_enable_valid(phi_dw_conv_s1_r_dw__x_013262_io_enable_valid),
    .io_enable_bits_control(phi_dw_conv_s1_r_dw__x_013262_io_enable_bits_control),
    .io_InData_0_ready(phi_dw_conv_s1_r_dw__x_013262_io_InData_0_ready),
    .io_InData_0_valid(phi_dw_conv_s1_r_dw__x_013262_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_dw_conv_s1_r_dw__x_013262_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi_dw_conv_s1_r_dw__x_013262_io_InData_1_ready),
    .io_InData_1_valid(phi_dw_conv_s1_r_dw__x_013262_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_dw_conv_s1_r_dw__x_013262_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_dw_conv_s1_r_dw__x_013262_io_InData_1_bits_data),
    .io_Mask_ready(phi_dw_conv_s1_r_dw__x_013262_io_Mask_ready),
    .io_Mask_valid(phi_dw_conv_s1_r_dw__x_013262_io_Mask_valid),
    .io_Mask_bits(phi_dw_conv_s1_r_dw__x_013262_io_Mask_bits),
    .io_Out_0_ready(phi_dw_conv_s1_r_dw__x_013262_io_Out_0_ready),
    .io_Out_0_valid(phi_dw_conv_s1_r_dw__x_013262_io_Out_0_valid),
    .io_Out_0_bits_data(phi_dw_conv_s1_r_dw__x_013262_io_Out_0_bits_data),
    .io_Out_1_ready(phi_dw_conv_s1_r_dw__x_013262_io_Out_1_ready),
    .io_Out_1_valid(phi_dw_conv_s1_r_dw__x_013262_io_Out_1_valid),
    .io_Out_1_bits_data(phi_dw_conv_s1_r_dw__x_013262_io_Out_1_bits_data)
  );
  ComputeNode_31 binaryOp_add3563 ( // @[extracted_function_reduction.scala 314:32]
    .clock(binaryOp_add3563_clock),
    .reset(binaryOp_add3563_reset),
    .io_enable_ready(binaryOp_add3563_io_enable_ready),
    .io_enable_valid(binaryOp_add3563_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add3563_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add3563_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add3563_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add3563_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add3563_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add3563_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add3563_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add3563_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add3563_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add3563_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add3563_io_RightIO_bits_data)
  );
  GepNode_1 Gep_arrayidx64 ( // @[extracted_function_reduction.scala 317:30]
    .clock(Gep_arrayidx64_clock),
    .reset(Gep_arrayidx64_reset),
    .io_enable_ready(Gep_arrayidx64_io_enable_ready),
    .io_enable_valid(Gep_arrayidx64_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx64_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx64_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx64_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx64_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx64_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx64_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx64_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx64_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx64_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx64_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx64_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx64_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx64_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx64_io_idx_0_bits_data)
  );
  UnTypLoad_1 ld_65 ( // @[extracted_function_reduction.scala 320:21]
    .clock(ld_65_clock),
    .reset(ld_65_reset),
    .io_enable_ready(ld_65_io_enable_ready),
    .io_enable_valid(ld_65_io_enable_valid),
    .io_enable_bits_taskID(ld_65_io_enable_bits_taskID),
    .io_enable_bits_control(ld_65_io_enable_bits_control),
    .io_Out_0_ready(ld_65_io_Out_0_ready),
    .io_Out_0_valid(ld_65_io_Out_0_valid),
    .io_Out_0_bits_data(ld_65_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_65_io_GepAddr_ready),
    .io_GepAddr_valid(ld_65_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_65_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_65_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_65_io_GepAddr_bits_data),
    .io_memReq_ready(ld_65_io_memReq_ready),
    .io_memReq_valid(ld_65_io_memReq_valid),
    .io_memReq_bits_address(ld_65_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_65_io_memReq_bits_taskID),
    .io_memResp_valid(ld_65_io_memResp_valid),
    .io_memResp_data(ld_65_io_memResp_data)
  );
  SextNode_1 sextconv3766 ( // @[extracted_function_reduction.scala 323:28]
    .clock(sextconv3766_clock),
    .reset(sextconv3766_reset),
    .io_Input_ready(sextconv3766_io_Input_ready),
    .io_Input_valid(sextconv3766_io_Input_valid),
    .io_Input_bits_data(sextconv3766_io_Input_bits_data),
    .io_enable_ready(sextconv3766_io_enable_ready),
    .io_enable_valid(sextconv3766_io_enable_valid),
    .io_enable_bits_taskID(sextconv3766_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv3766_io_Out_0_ready),
    .io_Out_0_valid(sextconv3766_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv3766_io_Out_0_bits_data)
  );
  ComputeNode_32 binaryOp_add3867 ( // @[extracted_function_reduction.scala 326:32]
    .clock(binaryOp_add3867_clock),
    .reset(binaryOp_add3867_reset),
    .io_enable_ready(binaryOp_add3867_io_enable_ready),
    .io_enable_valid(binaryOp_add3867_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add3867_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add3867_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add3867_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add3867_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add3867_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add3867_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add3867_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add3867_io_Out_1_valid),
    .io_Out_1_bits_taskID(binaryOp_add3867_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(binaryOp_add3867_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add3867_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add3867_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add3867_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add3867_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add3867_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add3867_io_RightIO_bits_data)
  );
  ComputeNode_33 binaryOp_inc68 ( // @[extracted_function_reduction.scala 329:30]
    .clock(binaryOp_inc68_clock),
    .reset(binaryOp_inc68_reset),
    .io_enable_ready(binaryOp_inc68_io_enable_ready),
    .io_enable_valid(binaryOp_inc68_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_inc68_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_inc68_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_inc68_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_inc68_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_inc68_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_inc68_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_inc68_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_inc68_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_inc68_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_inc68_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_inc68_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_inc68_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_inc68_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_inc68_io_RightIO_valid)
  );
  ComputeNode_34 icmp_exitcond69 ( // @[extracted_function_reduction.scala 332:31]
    .clock(icmp_exitcond69_clock),
    .reset(icmp_exitcond69_reset),
    .io_enable_ready(icmp_exitcond69_io_enable_ready),
    .io_enable_valid(icmp_exitcond69_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond69_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond69_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond69_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond69_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond69_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond69_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond69_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond69_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond69_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond69_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond69_io_RightIO_valid)
  );
  CBranchNodeVariable_8 br_70 ( // @[extracted_function_reduction.scala 335:21]
    .clock(br_70_clock),
    .reset(br_70_reset),
    .io_enable_ready(br_70_io_enable_ready),
    .io_enable_valid(br_70_io_enable_valid),
    .io_enable_bits_taskID(br_70_io_enable_bits_taskID),
    .io_enable_bits_control(br_70_io_enable_bits_control),
    .io_CmpIO_ready(br_70_io_CmpIO_ready),
    .io_CmpIO_valid(br_70_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_70_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_70_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_70_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_70_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_70_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_70_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_70_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_70_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_70_io_FalseOutput_0_bits_control)
  );
  ConstFastNode const0 ( // @[extracted_function_reduction.scala 344:22]
    .clock(const0_clock),
    .reset(const0_reset),
    .io_enable_ready(const0_io_enable_ready),
    .io_enable_valid(const0_io_enable_valid),
    .io_enable_bits_taskID(const0_io_enable_bits_taskID),
    .io_Out_ready(const0_io_Out_ready),
    .io_Out_valid(const0_io_Out_valid)
  );
  ConstFastNode_1 const1 ( // @[extracted_function_reduction.scala 347:22]
    .clock(const1_clock),
    .reset(const1_reset),
    .io_enable_ready(const1_io_enable_ready),
    .io_enable_valid(const1_io_enable_valid),
    .io_enable_bits_taskID(const1_io_enable_bits_taskID),
    .io_Out_ready(const1_io_Out_ready),
    .io_Out_valid(const1_io_Out_valid)
  );
  ConstFastNode_2 const2 ( // @[extracted_function_reduction.scala 350:22]
    .clock(const2_clock),
    .reset(const2_reset),
    .io_enable_ready(const2_io_enable_ready),
    .io_enable_valid(const2_io_enable_valid),
    .io_enable_bits_taskID(const2_io_enable_bits_taskID),
    .io_Out_ready(const2_io_Out_ready),
    .io_Out_valid(const2_io_Out_valid)
  );
  ConstFastNode_3 const3 ( // @[extracted_function_reduction.scala 353:22]
    .clock(const3_clock),
    .reset(const3_reset),
    .io_enable_ready(const3_io_enable_ready),
    .io_enable_valid(const3_io_enable_valid),
    .io_enable_bits_taskID(const3_io_enable_bits_taskID),
    .io_Out_ready(const3_io_Out_ready),
    .io_Out_valid(const3_io_Out_valid),
    .io_Out_bits_taskID(const3_io_Out_bits_taskID)
  );
  ConstFastNode_4 const4 ( // @[extracted_function_reduction.scala 356:22]
    .clock(const4_clock),
    .reset(const4_reset),
    .io_enable_ready(const4_io_enable_ready),
    .io_enable_valid(const4_io_enable_valid),
    .io_enable_bits_taskID(const4_io_enable_bits_taskID),
    .io_Out_ready(const4_io_Out_ready),
    .io_Out_valid(const4_io_Out_valid)
  );
  ConstFastNode_5 const5 ( // @[extracted_function_reduction.scala 359:22]
    .clock(const5_clock),
    .reset(const5_reset),
    .io_enable_ready(const5_io_enable_ready),
    .io_enable_valid(const5_io_enable_valid),
    .io_enable_bits_taskID(const5_io_enable_bits_taskID),
    .io_Out_ready(const5_io_Out_ready),
    .io_Out_valid(const5_io_Out_valid)
  );
  ConstFastNode_6 const6 ( // @[extracted_function_reduction.scala 362:22]
    .clock(const6_clock),
    .reset(const6_reset),
    .io_enable_ready(const6_io_enable_ready),
    .io_enable_valid(const6_io_enable_valid),
    .io_enable_bits_taskID(const6_io_enable_bits_taskID),
    .io_Out_ready(const6_io_Out_ready),
    .io_Out_valid(const6_io_Out_valid)
  );
  ConstFastNode_7 const7 ( // @[extracted_function_reduction.scala 365:22]
    .clock(const7_clock),
    .reset(const7_reset),
    .io_enable_ready(const7_io_enable_ready),
    .io_enable_valid(const7_io_enable_valid),
    .io_enable_bits_taskID(const7_io_enable_bits_taskID),
    .io_Out_ready(const7_io_Out_ready),
    .io_Out_valid(const7_io_Out_valid),
    .io_Out_bits_taskID(const7_io_Out_bits_taskID)
  );
  ConstFastNode_8 const8 ( // @[extracted_function_reduction.scala 368:22]
    .clock(const8_clock),
    .reset(const8_reset),
    .io_enable_ready(const8_io_enable_ready),
    .io_enable_valid(const8_io_enable_valid),
    .io_enable_bits_taskID(const8_io_enable_bits_taskID),
    .io_Out_ready(const8_io_Out_ready),
    .io_Out_valid(const8_io_Out_valid),
    .io_Out_bits_taskID(const8_io_Out_bits_taskID)
  );
  ConstFastNode_9 const9 ( // @[extracted_function_reduction.scala 371:22]
    .clock(const9_clock),
    .reset(const9_reset),
    .io_enable_ready(const9_io_enable_ready),
    .io_enable_valid(const9_io_enable_valid),
    .io_enable_bits_taskID(const9_io_enable_bits_taskID),
    .io_Out_ready(const9_io_Out_ready),
    .io_Out_valid(const9_io_Out_valid)
  );
  ConstFastNode_10 const10 ( // @[extracted_function_reduction.scala 374:23]
    .clock(const10_clock),
    .reset(const10_reset),
    .io_enable_ready(const10_io_enable_ready),
    .io_enable_valid(const10_io_enable_valid),
    .io_enable_bits_taskID(const10_io_enable_bits_taskID),
    .io_Out_ready(const10_io_Out_ready),
    .io_Out_valid(const10_io_Out_valid)
  );
  ConstFastNode_11 const11 ( // @[extracted_function_reduction.scala 377:23]
    .clock(const11_clock),
    .reset(const11_reset),
    .io_enable_ready(const11_io_enable_ready),
    .io_enable_valid(const11_io_enable_valid),
    .io_enable_bits_taskID(const11_io_enable_bits_taskID),
    .io_Out_ready(const11_io_Out_ready),
    .io_Out_valid(const11_io_Out_valid),
    .io_Out_bits_taskID(const11_io_Out_bits_taskID)
  );
  ConstFastNode_12 const12 ( // @[extracted_function_reduction.scala 380:23]
    .clock(const12_clock),
    .reset(const12_reset),
    .io_enable_ready(const12_io_enable_ready),
    .io_enable_valid(const12_io_enable_valid),
    .io_enable_bits_taskID(const12_io_enable_bits_taskID),
    .io_Out_ready(const12_io_Out_ready),
    .io_Out_valid(const12_io_Out_valid)
  );
  ConstFastNode_13 const13 ( // @[extracted_function_reduction.scala 383:23]
    .clock(const13_clock),
    .reset(const13_reset),
    .io_enable_ready(const13_io_enable_ready),
    .io_enable_valid(const13_io_enable_valid),
    .io_enable_bits_taskID(const13_io_enable_bits_taskID),
    .io_Out_ready(const13_io_Out_ready),
    .io_Out_valid(const13_io_Out_valid)
  );
  assign io_in_ready = InputSplitter_io_In_ready; // @[extracted_function_reduction.scala 54:23]
  assign io_MemReq_valid = MemCtrl_io_MemReq_valid; // @[extracted_function_reduction.scala 50:13]
  assign io_MemReq_bits_addr = MemCtrl_io_MemReq_bits_addr; // @[extracted_function_reduction.scala 50:13]
  assign io_MemReq_bits_data = MemCtrl_io_MemReq_bits_data; // @[extracted_function_reduction.scala 50:13]
  assign io_MemReq_bits_mask = MemCtrl_io_MemReq_bits_mask; // @[extracted_function_reduction.scala 50:13]
  assign io_MemReq_bits_tag = MemCtrl_io_MemReq_bits_tag; // @[extracted_function_reduction.scala 50:13]
  assign io_MemReq_bits_taskID = MemCtrl_io_MemReq_bits_taskID; // @[extracted_function_reduction.scala 50:13]
  assign io_MemReq_bits_iswrite = MemCtrl_io_MemReq_bits_iswrite; // @[extracted_function_reduction.scala 50:13]
  assign io_MemReq_bits_tile = 32'h0; // @[extracted_function_reduction.scala 50:13]
  assign io_out_valid = ret_9_io_Out_valid; // @[extracted_function_reduction.scala 1192:10]
  assign io_out_bits_enable_taskID = ret_9_io_Out_bits_enable_taskID; // @[extracted_function_reduction.scala 1192:10]
  assign io_out_bits_enable_control = ret_9_io_Out_bits_enable_control; // @[extracted_function_reduction.scala 1192:10]
  assign MemCtrl_clock = clock;
  assign MemCtrl_reset = reset;
  assign MemCtrl_io_WriteIn_0_valid = st_47_io_memReq_valid; // @[extracted_function_reduction.scala 1024:25]
  assign MemCtrl_io_WriteIn_0_bits_address = st_47_io_memReq_bits_address; // @[extracted_function_reduction.scala 1024:25]
  assign MemCtrl_io_WriteIn_0_bits_data = st_47_io_memReq_bits_data; // @[extracted_function_reduction.scala 1024:25]
  assign MemCtrl_io_WriteIn_0_bits_taskID = st_47_io_memReq_bits_taskID; // @[extracted_function_reduction.scala 1024:25]
  assign MemCtrl_io_ReadIn_0_valid = ld_45_io_memReq_valid; // @[extracted_function_reduction.scala 1020:24]
  assign MemCtrl_io_ReadIn_0_bits_address = ld_45_io_memReq_bits_address; // @[extracted_function_reduction.scala 1020:24]
  assign MemCtrl_io_ReadIn_0_bits_taskID = ld_45_io_memReq_bits_taskID; // @[extracted_function_reduction.scala 1020:24]
  assign MemCtrl_io_ReadIn_1_valid = ld_65_io_memReq_valid; // @[extracted_function_reduction.scala 1028:24]
  assign MemCtrl_io_ReadIn_1_bits_address = ld_65_io_memReq_bits_address; // @[extracted_function_reduction.scala 1028:24]
  assign MemCtrl_io_ReadIn_1_bits_taskID = ld_65_io_memReq_bits_taskID; // @[extracted_function_reduction.scala 1028:24]
  assign MemCtrl_io_MemResp_valid = io_MemResp_valid; // @[extracted_function_reduction.scala 51:22]
  assign MemCtrl_io_MemResp_bits_data = io_MemResp_bits_data; // @[extracted_function_reduction.scala 51:22]
  assign MemCtrl_io_MemResp_bits_tag = io_MemResp_bits_tag; // @[extracted_function_reduction.scala 51:22]
  assign MemCtrl_io_MemResp_bits_iswrite = io_MemResp_bits_iswrite; // @[extracted_function_reduction.scala 51:22]
  assign MemCtrl_io_MemReq_ready = io_MemReq_ready; // @[extracted_function_reduction.scala 50:13]
  assign InputSplitter_clock = clock;
  assign InputSplitter_reset = reset;
  assign InputSplitter_io_In_valid = io_in_valid; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_enable_taskID = io_in_bits_enable_taskID; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_enable_control = io_in_bits_enable_control; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field10_data = io_in_bits_data_field10_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field9_data = io_in_bits_data_field9_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field8_taskID = io_in_bits_data_field8_taskID; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field8_data = io_in_bits_data_field8_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field7_data = io_in_bits_data_field7_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field6_taskID = io_in_bits_data_field6_taskID; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field6_data = io_in_bits_data_field6_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field5_data = io_in_bits_data_field5_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field4_taskID = io_in_bits_data_field4_taskID; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field4_data = io_in_bits_data_field4_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field3_data = io_in_bits_data_field3_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field2_data = io_in_bits_data_field2_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field1_taskID = io_in_bits_data_field1_taskID; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field1_data = io_in_bits_data_field1_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field0_taskID = io_in_bits_data_field0_taskID; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_In_bits_data_field0_data = io_in_bits_data_field0_data; // @[extracted_function_reduction.scala 54:23]
  assign InputSplitter_io_Out_enable_ready = bb_entry0_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 391:31]
  assign InputSplitter_io_Out_data_field10_0_ready = Loop_5_io_InLiveIn_7_ready; // @[extracted_function_reduction.scala 595:25]
  assign InputSplitter_io_Out_data_field9_0_ready = binaryOp_add0_io_LeftIO_ready; // @[extracted_function_reduction.scala 1182:27]
  assign InputSplitter_io_Out_data_field8_0_ready = Loop_5_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 581:25]
  assign InputSplitter_io_Out_data_field8_1_ready = binaryOp_add0_io_RightIO_ready; // @[extracted_function_reduction.scala 1178:28]
  assign InputSplitter_io_Out_data_field8_2_ready = icmp_cmp1421_io_RightIO_ready; // @[extracted_function_reduction.scala 1180:27]
  assign InputSplitter_io_Out_data_field7_0_ready = Loop_5_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 583:25]
  assign InputSplitter_io_Out_data_field7_1_ready = binaryOp_add43_io_LeftIO_ready; // @[extracted_function_reduction.scala 1176:28]
  assign InputSplitter_io_Out_data_field6_0_ready = Loop_5_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 587:25]
  assign InputSplitter_io_Out_data_field6_1_ready = binaryOp_add43_io_RightIO_ready; // @[extracted_function_reduction.scala 1172:29]
  assign InputSplitter_io_Out_data_field6_2_ready = icmp_cmp51394_io_RightIO_ready; // @[extracted_function_reduction.scala 1174:28]
  assign InputSplitter_io_Out_data_field5_0_ready = Loop_5_io_InLiveIn_5_ready; // @[extracted_function_reduction.scala 591:25]
  assign InputSplitter_io_Out_data_field5_1_ready = binaryOp_add125_io_LeftIO_ready; // @[extracted_function_reduction.scala 1170:29]
  assign InputSplitter_io_Out_data_field4_0_ready = Loop_5_io_InLiveIn_6_ready; // @[extracted_function_reduction.scala 593:25]
  assign InputSplitter_io_Out_data_field4_1_ready = binaryOp_add125_io_RightIO_ready; // @[extracted_function_reduction.scala 1166:30]
  assign InputSplitter_io_Out_data_field4_2_ready = icmp_cmp131376_io_RightIO_ready; // @[extracted_function_reduction.scala 1168:29]
  assign InputSplitter_io_Out_data_field3_0_ready = Loop_5_io_InLiveIn_9_ready; // @[extracted_function_reduction.scala 599:25]
  assign InputSplitter_io_Out_data_field2_0_ready = Loop_5_io_InLiveIn_10_ready; // @[extracted_function_reduction.scala 601:26]
  assign InputSplitter_io_Out_data_field1_0_ready = Loop_5_io_InLiveIn_11_ready; // @[extracted_function_reduction.scala 603:26]
  assign InputSplitter_io_Out_data_field0_0_ready = Loop_5_io_InLiveIn_8_ready; // @[extracted_function_reduction.scala 597:25]
  assign Loop_0_clock = clock;
  assign Loop_0_reset = reset;
  assign Loop_0_io_enable_valid = br_56_io_Out_0_valid; // @[extracted_function_reduction.scala 465:20]
  assign Loop_0_io_enable_bits_taskID = br_56_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 465:20]
  assign Loop_0_io_enable_bits_control = br_56_io_Out_0_bits_control; // @[extracted_function_reduction.scala 465:20]
  assign Loop_0_io_InLiveIn_0_valid = phi_dw_conv_013551_io_Out_0_valid; // @[extracted_function_reduction.scala 513:25]
  assign Loop_0_io_InLiveIn_0_bits_taskID = phi_dw_conv_013551_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 513:25]
  assign Loop_0_io_InLiveIn_0_bits_data = phi_dw_conv_013551_io_Out_0_bits_data; // @[extracted_function_reduction.scala 513:25]
  assign Loop_0_io_InLiveIn_1_valid = binaryOp_add3055_io_Out_0_valid; // @[extracted_function_reduction.scala 515:25]
  assign Loop_0_io_InLiveIn_1_bits_data = binaryOp_add3055_io_Out_0_bits_data; // @[extracted_function_reduction.scala 515:25]
  assign Loop_0_io_InLiveIn_2_valid = Loop_1_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 517:25]
  assign Loop_0_io_InLiveIn_2_bits_taskID = Loop_1_io_OutLiveIn_field1_0_bits_taskID; // @[extracted_function_reduction.scala 517:25]
  assign Loop_0_io_InLiveIn_2_bits_data = Loop_1_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 517:25]
  assign Loop_0_io_OutLiveIn_field2_0_ready = Gep_arrayidx64_io_baseAddress_ready; // @[extracted_function_reduction.scala 621:33]
  assign Loop_0_io_OutLiveIn_field1_0_ready = binaryOp_add3563_io_LeftIO_ready; // @[extracted_function_reduction.scala 619:30]
  assign Loop_0_io_OutLiveIn_field0_0_ready = phi_dw_conv_113361_io_InData_0_ready; // @[extracted_function_reduction.scala 617:35]
  assign Loop_0_io_activate_loop_start_ready = bb_for_body3418_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 449:37]
  assign Loop_0_io_activate_loop_back_ready = bb_for_body3418_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 451:37]
  assign Loop_0_io_loopBack_0_valid = br_70_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 467:25]
  assign Loop_0_io_loopBack_0_bits_taskID = br_70_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 467:25]
  assign Loop_0_io_loopBack_0_bits_control = br_70_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 467:25]
  assign Loop_0_io_loopFinish_0_valid = br_70_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 469:27]
  assign Loop_0_io_loopFinish_0_bits_control = br_70_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 469:27]
  assign Loop_0_io_CarryDepenIn_0_valid = binaryOp_add3867_io_Out_1_valid; // @[extracted_function_reduction.scala 697:29]
  assign Loop_0_io_CarryDepenIn_0_bits_taskID = binaryOp_add3867_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 697:29]
  assign Loop_0_io_CarryDepenIn_0_bits_data = binaryOp_add3867_io_Out_1_bits_data; // @[extracted_function_reduction.scala 697:29]
  assign Loop_0_io_CarryDepenIn_1_valid = binaryOp_inc68_io_Out_0_valid; // @[extracted_function_reduction.scala 699:29]
  assign Loop_0_io_CarryDepenIn_1_bits_taskID = binaryOp_inc68_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 699:29]
  assign Loop_0_io_CarryDepenIn_1_bits_data = binaryOp_inc68_io_Out_0_bits_data; // @[extracted_function_reduction.scala 699:29]
  assign Loop_0_io_CarryDepenOut_field1_0_ready = phi_dw_conv_s1_r_dw__x_013262_io_InData_1_ready; // @[extracted_function_reduction.scala 721:46]
  assign Loop_0_io_CarryDepenOut_field0_0_ready = phi_dw_conv_113361_io_InData_1_ready; // @[extracted_function_reduction.scala 719:35]
  assign Loop_0_io_InLiveOut_0_valid = binaryOp_add3867_io_Out_0_valid; // @[extracted_function_reduction.scala 677:26]
  assign Loop_0_io_InLiveOut_0_bits_taskID = binaryOp_add3867_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 677:26]
  assign Loop_0_io_InLiveOut_0_bits_data = binaryOp_add3867_io_Out_0_bits_data; // @[extracted_function_reduction.scala 677:26]
  assign Loop_0_io_OutLiveOut_field0_0_ready = phiadd38_lcssa57_io_InData_0_ready; // @[extracted_function_reduction.scala 687:33]
  assign Loop_0_io_loopExit_0_ready = bb_for_cond_cleanup3317_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 447:45]
  assign Loop_1_clock = clock;
  assign Loop_1_reset = reset;
  assign Loop_1_io_enable_valid = br_41_io_Out_0_valid; // @[extracted_function_reduction.scala 471:20]
  assign Loop_1_io_enable_bits_taskID = br_41_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 471:20]
  assign Loop_1_io_enable_bits_control = br_41_io_Out_0_bits_control; // @[extracted_function_reduction.scala 471:20]
  assign Loop_1_io_InLiveIn_0_valid = binaryOp_add2340_io_Out_0_valid; // @[extracted_function_reduction.scala 519:25]
  assign Loop_1_io_InLiveIn_0_bits_data = binaryOp_add2340_io_Out_0_bits_data; // @[extracted_function_reduction.scala 519:25]
  assign Loop_1_io_InLiveIn_1_valid = Loop_2_io_OutLiveIn_field4_0_valid; // @[extracted_function_reduction.scala 521:25]
  assign Loop_1_io_InLiveIn_1_bits_taskID = Loop_2_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_reduction.scala 521:25]
  assign Loop_1_io_InLiveIn_1_bits_data = Loop_2_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_reduction.scala 521:25]
  assign Loop_1_io_InLiveIn_2_valid = Loop_2_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 523:25]
  assign Loop_1_io_InLiveIn_2_bits_data = Loop_2_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 523:25]
  assign Loop_1_io_InLiveIn_3_valid = Loop_2_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 525:25]
  assign Loop_1_io_InLiveIn_3_bits_data = Loop_2_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 525:25]
  assign Loop_1_io_OutLiveIn_field3_0_ready = binaryOp_add2853_io_RightIO_ready; // @[extracted_function_reduction.scala 627:31]
  assign Loop_1_io_OutLiveIn_field2_0_ready = binaryOp_mul2954_io_RightIO_ready; // @[extracted_function_reduction.scala 625:31]
  assign Loop_1_io_OutLiveIn_field1_0_ready = Loop_0_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 517:25]
  assign Loop_1_io_OutLiveIn_field0_0_ready = binaryOp_add3055_io_LeftIO_ready; // @[extracted_function_reduction.scala 623:30]
  assign Loop_1_io_activate_loop_start_ready = bb_for_body2716_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 443:37]
  assign Loop_1_io_activate_loop_back_ready = bb_for_body2716_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 445:37]
  assign Loop_1_io_loopBack_0_valid = br_60_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 473:25]
  assign Loop_1_io_loopBack_0_bits_taskID = br_60_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 473:25]
  assign Loop_1_io_loopBack_0_bits_control = br_60_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 473:25]
  assign Loop_1_io_loopFinish_0_valid = br_60_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 475:27]
  assign Loop_1_io_loopFinish_0_bits_control = br_60_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 475:27]
  assign Loop_1_io_CarryDepenIn_0_valid = binaryOp_inc4158_io_Out_0_valid; // @[extracted_function_reduction.scala 701:29]
  assign Loop_1_io_CarryDepenIn_0_bits_taskID = binaryOp_inc4158_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 701:29]
  assign Loop_1_io_CarryDepenIn_0_bits_data = binaryOp_inc4158_io_Out_0_bits_data; // @[extracted_function_reduction.scala 701:29]
  assign Loop_1_io_CarryDepenIn_1_valid = phiadd38_lcssa57_io_Out_1_valid; // @[extracted_function_reduction.scala 703:29]
  assign Loop_1_io_CarryDepenIn_1_bits_taskID = phiadd38_lcssa57_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 703:29]
  assign Loop_1_io_CarryDepenIn_1_bits_data = phiadd38_lcssa57_io_Out_1_bits_data; // @[extracted_function_reduction.scala 703:29]
  assign Loop_1_io_CarryDepenOut_field1_0_ready = phi_dw_conv_013551_io_InData_1_ready; // @[extracted_function_reduction.scala 725:35]
  assign Loop_1_io_CarryDepenOut_field0_0_ready = phi_dw_conv_s1_r_dw__y_013452_io_InData_1_ready; // @[extracted_function_reduction.scala 723:46]
  assign Loop_1_io_InLiveOut_0_valid = phiadd38_lcssa57_io_Out_0_valid; // @[extracted_function_reduction.scala 679:26]
  assign Loop_1_io_InLiveOut_0_bits_taskID = phiadd38_lcssa57_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 679:26]
  assign Loop_1_io_InLiveOut_0_bits_data = phiadd38_lcssa57_io_Out_0_bits_data; // @[extracted_function_reduction.scala 679:26]
  assign Loop_1_io_OutLiveOut_field0_0_ready = phiadd38_lcssa_lcssa42_io_InData_0_ready; // @[extracted_function_reduction.scala 689:39]
  assign Loop_1_io_loopExit_0_ready = bb_for_cond_cleanup2615_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 441:45]
  assign Loop_2_clock = clock;
  assign Loop_2_reset = reset;
  assign Loop_2_io_enable_valid = br_34_io_Out_0_valid; // @[extracted_function_reduction.scala 477:20]
  assign Loop_2_io_enable_bits_taskID = br_34_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 477:20]
  assign Loop_2_io_enable_bits_control = br_34_io_Out_0_bits_control; // @[extracted_function_reduction.scala 477:20]
  assign Loop_2_io_InLiveIn_0_valid = binaryOp_sub1630_io_Out_0_valid; // @[extracted_function_reduction.scala 527:25]
  assign Loop_2_io_InLiveIn_0_bits_data = binaryOp_sub1630_io_Out_0_bits_data; // @[extracted_function_reduction.scala 527:25]
  assign Loop_2_io_InLiveIn_1_valid = Gep_arrayidx5033_io_Out_0_valid; // @[extracted_function_reduction.scala 529:25]
  assign Loop_2_io_InLiveIn_1_bits_predicate = Gep_arrayidx5033_io_Out_0_bits_predicate; // @[extracted_function_reduction.scala 529:25]
  assign Loop_2_io_InLiveIn_1_bits_taskID = Gep_arrayidx5033_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 529:25]
  assign Loop_2_io_InLiveIn_1_bits_data = Gep_arrayidx5033_io_Out_0_bits_data; // @[extracted_function_reduction.scala 529:25]
  assign Loop_2_io_InLiveIn_2_valid = Loop_3_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 531:25]
  assign Loop_2_io_InLiveIn_2_bits_data = Loop_3_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 531:25]
  assign Loop_2_io_InLiveIn_3_valid = Loop_3_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 533:25]
  assign Loop_2_io_InLiveIn_3_bits_data = Loop_3_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 533:25]
  assign Loop_2_io_InLiveIn_4_valid = Loop_3_io_OutLiveIn_field4_0_valid; // @[extracted_function_reduction.scala 535:25]
  assign Loop_2_io_InLiveIn_4_bits_taskID = Loop_3_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_reduction.scala 535:25]
  assign Loop_2_io_InLiveIn_4_bits_data = Loop_3_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_reduction.scala 535:25]
  assign Loop_2_io_InLiveIn_5_valid = Loop_3_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 537:25]
  assign Loop_2_io_InLiveIn_5_bits_data = Loop_3_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 537:25]
  assign Loop_2_io_OutLiveIn_field5_0_ready = binaryOp_mul2239_io_RightIO_ready; // @[extracted_function_reduction.scala 635:31]
  assign Loop_2_io_OutLiveIn_field4_0_ready = Loop_1_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 521:25]
  assign Loop_2_io_OutLiveIn_field3_0_ready = Loop_1_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 525:25]
  assign Loop_2_io_OutLiveIn_field2_0_ready = Loop_1_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 523:25]
  assign Loop_2_io_OutLiveIn_field1_0_ready = ld_45_io_GepAddr_ready; // @[extracted_function_reduction.scala 631:20]
  assign Loop_2_io_OutLiveIn_field1_1_ready = st_47_io_GepAddr_ready; // @[extracted_function_reduction.scala 633:20]
  assign Loop_2_io_OutLiveIn_field0_0_ready = binaryOp_add2340_io_LeftIO_ready; // @[extracted_function_reduction.scala 629:30]
  assign Loop_2_io_activate_loop_start_ready = bb_for_body2114_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 437:37]
  assign Loop_2_io_activate_loop_back_ready = bb_for_body2114_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 439:37]
  assign Loop_2_io_loopBack_0_valid = br_50_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 479:25]
  assign Loop_2_io_loopBack_0_bits_taskID = br_50_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 479:25]
  assign Loop_2_io_loopBack_0_bits_control = br_50_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 479:25]
  assign Loop_2_io_loopFinish_0_valid = br_50_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 481:27]
  assign Loop_2_io_loopFinish_0_bits_control = br_50_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 481:27]
  assign Loop_2_io_CarryDepenIn_0_valid = binaryOp_inc5548_io_Out_0_valid; // @[extracted_function_reduction.scala 705:29]
  assign Loop_2_io_CarryDepenIn_0_bits_taskID = binaryOp_inc5548_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 705:29]
  assign Loop_2_io_CarryDepenIn_0_bits_data = binaryOp_inc5548_io_Out_0_bits_data; // @[extracted_function_reduction.scala 705:29]
  assign Loop_2_io_CarryDepenOut_field0_0_ready = phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_ready; // @[extracted_function_reduction.scala 727:56]
  assign Loop_2_io_loopExit_0_ready = bb_for_cond_cleanup2013_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 435:45]
  assign Loop_3_clock = clock;
  assign Loop_3_reset = reset;
  assign Loop_3_io_enable_valid = br_24_io_Out_0_valid; // @[extracted_function_reduction.scala 483:20]
  assign Loop_3_io_enable_bits_taskID = br_24_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 483:20]
  assign Loop_3_io_enable_bits_control = br_24_io_Out_0_bits_control; // @[extracted_function_reduction.scala 483:20]
  assign Loop_3_io_InLiveIn_0_valid = binaryOp_reass_mul23_io_Out_0_valid; // @[extracted_function_reduction.scala 539:25]
  assign Loop_3_io_InLiveIn_0_bits_data = binaryOp_reass_mul23_io_Out_0_bits_data; // @[extracted_function_reduction.scala 539:25]
  assign Loop_3_io_InLiveIn_1_valid = phi_pw_conv_reduction_s1_y_014019_io_Out_0_valid; // @[extracted_function_reduction.scala 541:25]
  assign Loop_3_io_InLiveIn_1_bits_data = phi_pw_conv_reduction_s1_y_014019_io_Out_0_bits_data; // @[extracted_function_reduction.scala 541:25]
  assign Loop_3_io_InLiveIn_2_valid = Loop_4_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 543:25]
  assign Loop_3_io_InLiveIn_2_bits_data = Loop_4_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 543:25]
  assign Loop_3_io_InLiveIn_3_valid = Loop_4_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 545:25]
  assign Loop_3_io_InLiveIn_3_bits_data = Loop_4_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 545:25]
  assign Loop_3_io_InLiveIn_4_valid = Loop_4_io_OutLiveIn_field4_0_valid; // @[extracted_function_reduction.scala 547:25]
  assign Loop_3_io_InLiveIn_4_bits_taskID = Loop_4_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_reduction.scala 547:25]
  assign Loop_3_io_InLiveIn_4_bits_data = Loop_4_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_reduction.scala 547:25]
  assign Loop_3_io_InLiveIn_5_valid = Loop_4_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 549:25]
  assign Loop_3_io_InLiveIn_5_bits_taskID = Loop_4_io_OutLiveIn_field3_0_bits_taskID; // @[extracted_function_reduction.scala 549:25]
  assign Loop_3_io_InLiveIn_5_bits_data = Loop_4_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 549:25]
  assign Loop_3_io_InLiveIn_6_valid = Loop_4_io_OutLiveIn_field5_0_valid; // @[extracted_function_reduction.scala 551:25]
  assign Loop_3_io_InLiveIn_6_bits_data = Loop_4_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_reduction.scala 551:25]
  assign Loop_3_io_InLiveIn_7_valid = Loop_4_io_OutLiveIn_field6_0_valid; // @[extracted_function_reduction.scala 553:25]
  assign Loop_3_io_InLiveIn_7_bits_data = Loop_4_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_reduction.scala 553:25]
  assign Loop_3_io_InLiveIn_8_valid = Loop_4_io_OutLiveIn_field7_0_valid; // @[extracted_function_reduction.scala 555:25]
  assign Loop_3_io_InLiveIn_8_bits_taskID = Loop_4_io_OutLiveIn_field7_0_bits_taskID; // @[extracted_function_reduction.scala 555:25]
  assign Loop_3_io_InLiveIn_8_bits_data = Loop_4_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_reduction.scala 555:25]
  assign Loop_3_io_OutLiveIn_field8_0_ready = phi_pw_conv_reduction_s1_x_013829_io_InData_0_ready; // @[extracted_function_reduction.scala 645:50]
  assign Loop_3_io_OutLiveIn_field8_1_ready = binaryOp_add1031_io_RightIO_ready; // @[extracted_function_reduction.scala 647:31]
  assign Loop_3_io_OutLiveIn_field7_0_ready = binaryOp_sub1630_io_RightIO_ready; // @[extracted_function_reduction.scala 643:31]
  assign Loop_3_io_OutLiveIn_field6_0_ready = icmp_exitcond14636_io_RightIO_ready; // @[extracted_function_reduction.scala 641:33]
  assign Loop_3_io_OutLiveIn_field5_0_ready = Gep_arrayidx5033_io_baseAddress_ready; // @[extracted_function_reduction.scala 639:35]
  assign Loop_3_io_OutLiveIn_field4_0_ready = Loop_2_io_InLiveIn_4_ready; // @[extracted_function_reduction.scala 535:25]
  assign Loop_3_io_OutLiveIn_field3_0_ready = Loop_2_io_InLiveIn_5_ready; // @[extracted_function_reduction.scala 537:25]
  assign Loop_3_io_OutLiveIn_field2_0_ready = Loop_2_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 531:25]
  assign Loop_3_io_OutLiveIn_field1_0_ready = Loop_2_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 533:25]
  assign Loop_3_io_OutLiveIn_field0_0_ready = binaryOp_add1732_io_RightIO_ready; // @[extracted_function_reduction.scala 637:31]
  assign Loop_3_io_activate_loop_start_ready = bb_for_body1512_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 431:37]
  assign Loop_3_io_activate_loop_back_ready = bb_for_body1512_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 433:37]
  assign Loop_3_io_loopBack_0_valid = br_37_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 485:25]
  assign Loop_3_io_loopBack_0_bits_taskID = br_37_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 485:25]
  assign Loop_3_io_loopBack_0_bits_control = br_37_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 485:25]
  assign Loop_3_io_loopFinish_0_valid = br_37_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 487:27]
  assign Loop_3_io_loopFinish_0_bits_control = br_37_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 487:27]
  assign Loop_3_io_CarryDepenIn_0_valid = binaryOp_inc5835_io_Out_0_valid; // @[extracted_function_reduction.scala 707:29]
  assign Loop_3_io_CarryDepenIn_0_bits_taskID = binaryOp_inc5835_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 707:29]
  assign Loop_3_io_CarryDepenIn_0_bits_data = binaryOp_inc5835_io_Out_0_bits_data; // @[extracted_function_reduction.scala 707:29]
  assign Loop_3_io_CarryDepenOut_field0_0_ready = phi_pw_conv_reduction_s1_x_013829_io_InData_1_ready; // @[extracted_function_reduction.scala 729:50]
  assign Loop_3_io_loopExit_0_ready = bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 429:54]
  assign Loop_4_clock = clock;
  assign Loop_4_reset = reset;
  assign Loop_4_io_enable_valid = br_14_io_Out_0_valid; // @[extracted_function_reduction.scala 489:20]
  assign Loop_4_io_enable_bits_taskID = br_14_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 489:20]
  assign Loop_4_io_enable_bits_control = br_14_io_Out_0_bits_control; // @[extracted_function_reduction.scala 489:20]
  assign Loop_4_io_InLiveIn_0_valid = binaryOp_mul112_io_Out_0_valid; // @[extracted_function_reduction.scala 557:25]
  assign Loop_4_io_InLiveIn_0_bits_data = binaryOp_mul112_io_Out_0_bits_data; // @[extracted_function_reduction.scala 557:25]
  assign Loop_4_io_InLiveIn_1_valid = Loop_5_io_OutLiveIn_field10_0_valid; // @[extracted_function_reduction.scala 559:25]
  assign Loop_4_io_InLiveIn_1_bits_data = Loop_5_io_OutLiveIn_field10_0_bits_data; // @[extracted_function_reduction.scala 559:25]
  assign Loop_4_io_InLiveIn_2_valid = Loop_5_io_OutLiveIn_field9_0_valid; // @[extracted_function_reduction.scala 561:25]
  assign Loop_4_io_InLiveIn_2_bits_data = Loop_5_io_OutLiveIn_field9_0_bits_data; // @[extracted_function_reduction.scala 561:25]
  assign Loop_4_io_InLiveIn_3_valid = Loop_5_io_OutLiveIn_field8_0_valid; // @[extracted_function_reduction.scala 563:25]
  assign Loop_4_io_InLiveIn_3_bits_taskID = Loop_5_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_reduction.scala 563:25]
  assign Loop_4_io_InLiveIn_3_bits_data = Loop_5_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_reduction.scala 563:25]
  assign Loop_4_io_InLiveIn_4_valid = Loop_5_io_OutLiveIn_field11_0_valid; // @[extracted_function_reduction.scala 565:25]
  assign Loop_4_io_InLiveIn_4_bits_taskID = Loop_5_io_OutLiveIn_field11_0_bits_taskID; // @[extracted_function_reduction.scala 565:25]
  assign Loop_4_io_InLiveIn_4_bits_data = Loop_5_io_OutLiveIn_field11_0_bits_data; // @[extracted_function_reduction.scala 565:25]
  assign Loop_4_io_InLiveIn_5_valid = Loop_5_io_OutLiveIn_field12_0_valid; // @[extracted_function_reduction.scala 567:25]
  assign Loop_4_io_InLiveIn_5_bits_data = Loop_5_io_OutLiveIn_field12_0_bits_data; // @[extracted_function_reduction.scala 567:25]
  assign Loop_4_io_InLiveIn_6_valid = Loop_5_io_OutLiveIn_field7_0_valid; // @[extracted_function_reduction.scala 569:25]
  assign Loop_4_io_InLiveIn_6_bits_data = Loop_5_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_reduction.scala 569:25]
  assign Loop_4_io_InLiveIn_7_valid = Loop_5_io_OutLiveIn_field6_0_valid; // @[extracted_function_reduction.scala 571:25]
  assign Loop_4_io_InLiveIn_7_bits_taskID = Loop_5_io_OutLiveIn_field6_0_bits_taskID; // @[extracted_function_reduction.scala 571:25]
  assign Loop_4_io_InLiveIn_7_bits_data = Loop_5_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_reduction.scala 571:25]
  assign Loop_4_io_InLiveIn_8_valid = Loop_5_io_OutLiveIn_field4_0_valid; // @[extracted_function_reduction.scala 573:25]
  assign Loop_4_io_InLiveIn_8_bits_taskID = Loop_5_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_reduction.scala 573:25]
  assign Loop_4_io_InLiveIn_8_bits_data = Loop_5_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_reduction.scala 573:25]
  assign Loop_4_io_InLiveIn_9_valid = Loop_5_io_OutLiveIn_field13_0_valid; // @[extracted_function_reduction.scala 575:25]
  assign Loop_4_io_InLiveIn_9_bits_data = Loop_5_io_OutLiveIn_field13_0_bits_data; // @[extracted_function_reduction.scala 575:25]
  assign Loop_4_io_InLiveIn_10_valid = Loop_5_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 577:26]
  assign Loop_4_io_InLiveIn_10_bits_taskID = Loop_5_io_OutLiveIn_field3_0_bits_taskID; // @[extracted_function_reduction.scala 577:26]
  assign Loop_4_io_InLiveIn_10_bits_data = Loop_5_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 577:26]
  assign Loop_4_io_InLiveIn_11_valid = Loop_5_io_OutLiveIn_field5_0_valid; // @[extracted_function_reduction.scala 579:26]
  assign Loop_4_io_InLiveIn_11_bits_data = Loop_5_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_reduction.scala 579:26]
  assign Loop_4_io_OutLiveIn_field11_0_ready = binaryOp_reass_mul23_io_RightIO_ready; // @[extracted_function_reduction.scala 659:35]
  assign Loop_4_io_OutLiveIn_field10_0_ready = phi_pw_conv_reduction_s1_y_014019_io_InData_1_ready; // @[extracted_function_reduction.scala 655:50]
  assign Loop_4_io_OutLiveIn_field10_1_ready = binaryOp_sub821_io_RightIO_ready; // @[extracted_function_reduction.scala 657:30]
  assign Loop_4_io_OutLiveIn_field9_0_ready = icmp_exitcond14727_io_RightIO_ready; // @[extracted_function_reduction.scala 653:33]
  assign Loop_4_io_OutLiveIn_field8_0_ready = br_20_io_CmpIO_ready; // @[extracted_function_reduction.scala 651:18]
  assign Loop_4_io_OutLiveIn_field7_0_ready = Loop_3_io_InLiveIn_8_ready; // @[extracted_function_reduction.scala 555:25]
  assign Loop_4_io_OutLiveIn_field6_0_ready = Loop_3_io_InLiveIn_7_ready; // @[extracted_function_reduction.scala 553:25]
  assign Loop_4_io_OutLiveIn_field5_0_ready = Loop_3_io_InLiveIn_6_ready; // @[extracted_function_reduction.scala 551:25]
  assign Loop_4_io_OutLiveIn_field4_0_ready = Loop_3_io_InLiveIn_4_ready; // @[extracted_function_reduction.scala 547:25]
  assign Loop_4_io_OutLiveIn_field3_0_ready = Loop_3_io_InLiveIn_5_ready; // @[extracted_function_reduction.scala 549:25]
  assign Loop_4_io_OutLiveIn_field2_0_ready = Loop_3_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 545:25]
  assign Loop_4_io_OutLiveIn_field1_0_ready = Loop_3_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 543:25]
  assign Loop_4_io_OutLiveIn_field0_0_ready = binaryOp_reass_add22_io_RightIO_ready; // @[extracted_function_reduction.scala 649:35]
  assign Loop_4_io_activate_loop_start_ready = bb_for_body78_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 425:35]
  assign Loop_4_io_activate_loop_back_ready = bb_for_body78_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 427:35]
  assign Loop_4_io_loopBack_0_valid = br_28_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 491:25]
  assign Loop_4_io_loopBack_0_bits_taskID = br_28_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 491:25]
  assign Loop_4_io_loopBack_0_bits_control = br_28_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 491:25]
  assign Loop_4_io_loopFinish_0_valid = br_28_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 493:27]
  assign Loop_4_io_loopFinish_0_bits_control = br_28_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 493:27]
  assign Loop_4_io_CarryDepenIn_0_valid = binaryOp_inc6126_io_Out_0_valid; // @[extracted_function_reduction.scala 709:29]
  assign Loop_4_io_CarryDepenIn_0_bits_taskID = binaryOp_inc6126_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 709:29]
  assign Loop_4_io_CarryDepenIn_0_bits_data = binaryOp_inc6126_io_Out_0_bits_data; // @[extracted_function_reduction.scala 709:29]
  assign Loop_4_io_CarryDepenOut_field0_0_ready = phi_pw_conv_reduction_s1_y_014019_io_InData_0_ready; // @[extracted_function_reduction.scala 731:50]
  assign Loop_4_io_loopExit_0_ready = bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 423:52]
  assign Loop_5_clock = clock;
  assign Loop_5_reset = reset;
  assign Loop_5_io_enable_valid = br_7_io_Out_0_valid; // @[extracted_function_reduction.scala 495:20]
  assign Loop_5_io_enable_bits_taskID = br_7_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 495:20]
  assign Loop_5_io_enable_bits_control = br_7_io_Out_0_bits_control; // @[extracted_function_reduction.scala 495:20]
  assign Loop_5_io_InLiveIn_0_valid = InputSplitter_io_Out_data_field8_0_valid; // @[extracted_function_reduction.scala 581:25]
  assign Loop_5_io_InLiveIn_0_bits_taskID = InputSplitter_io_Out_data_field8_0_bits_taskID; // @[extracted_function_reduction.scala 581:25]
  assign Loop_5_io_InLiveIn_0_bits_data = InputSplitter_io_Out_data_field8_0_bits_data; // @[extracted_function_reduction.scala 581:25]
  assign Loop_5_io_InLiveIn_1_valid = InputSplitter_io_Out_data_field7_0_valid; // @[extracted_function_reduction.scala 583:25]
  assign Loop_5_io_InLiveIn_1_bits_data = InputSplitter_io_Out_data_field7_0_bits_data; // @[extracted_function_reduction.scala 583:25]
  assign Loop_5_io_InLiveIn_2_valid = icmp_cmp51394_io_Out_0_valid; // @[extracted_function_reduction.scala 585:25]
  assign Loop_5_io_InLiveIn_2_bits_taskID = icmp_cmp51394_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 585:25]
  assign Loop_5_io_InLiveIn_2_bits_data = icmp_cmp51394_io_Out_0_bits_data; // @[extracted_function_reduction.scala 585:25]
  assign Loop_5_io_InLiveIn_3_valid = InputSplitter_io_Out_data_field6_0_valid; // @[extracted_function_reduction.scala 587:25]
  assign Loop_5_io_InLiveIn_3_bits_taskID = InputSplitter_io_Out_data_field6_0_bits_taskID; // @[extracted_function_reduction.scala 587:25]
  assign Loop_5_io_InLiveIn_3_bits_data = InputSplitter_io_Out_data_field6_0_bits_data; // @[extracted_function_reduction.scala 587:25]
  assign Loop_5_io_InLiveIn_4_valid = icmp_cmp131376_io_Out_0_valid; // @[extracted_function_reduction.scala 589:25]
  assign Loop_5_io_InLiveIn_4_bits_taskID = icmp_cmp131376_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 589:25]
  assign Loop_5_io_InLiveIn_4_bits_data = icmp_cmp131376_io_Out_0_bits_data; // @[extracted_function_reduction.scala 589:25]
  assign Loop_5_io_InLiveIn_5_valid = InputSplitter_io_Out_data_field5_0_valid; // @[extracted_function_reduction.scala 591:25]
  assign Loop_5_io_InLiveIn_5_bits_data = InputSplitter_io_Out_data_field5_0_bits_data; // @[extracted_function_reduction.scala 591:25]
  assign Loop_5_io_InLiveIn_6_valid = InputSplitter_io_Out_data_field4_0_valid; // @[extracted_function_reduction.scala 593:25]
  assign Loop_5_io_InLiveIn_6_bits_taskID = InputSplitter_io_Out_data_field4_0_bits_taskID; // @[extracted_function_reduction.scala 593:25]
  assign Loop_5_io_InLiveIn_6_bits_data = InputSplitter_io_Out_data_field4_0_bits_data; // @[extracted_function_reduction.scala 593:25]
  assign Loop_5_io_InLiveIn_7_valid = InputSplitter_io_Out_data_field10_0_valid; // @[extracted_function_reduction.scala 595:25]
  assign Loop_5_io_InLiveIn_7_bits_data = InputSplitter_io_Out_data_field10_0_bits_data; // @[extracted_function_reduction.scala 595:25]
  assign Loop_5_io_InLiveIn_8_valid = InputSplitter_io_Out_data_field0_0_valid; // @[extracted_function_reduction.scala 597:25]
  assign Loop_5_io_InLiveIn_8_bits_taskID = InputSplitter_io_Out_data_field0_0_bits_taskID; // @[extracted_function_reduction.scala 597:25]
  assign Loop_5_io_InLiveIn_8_bits_data = InputSplitter_io_Out_data_field0_0_bits_data; // @[extracted_function_reduction.scala 597:25]
  assign Loop_5_io_InLiveIn_9_valid = InputSplitter_io_Out_data_field3_0_valid; // @[extracted_function_reduction.scala 599:25]
  assign Loop_5_io_InLiveIn_9_bits_data = InputSplitter_io_Out_data_field3_0_bits_data; // @[extracted_function_reduction.scala 599:25]
  assign Loop_5_io_InLiveIn_10_valid = InputSplitter_io_Out_data_field2_0_valid; // @[extracted_function_reduction.scala 601:26]
  assign Loop_5_io_InLiveIn_10_bits_data = InputSplitter_io_Out_data_field2_0_bits_data; // @[extracted_function_reduction.scala 601:26]
  assign Loop_5_io_InLiveIn_11_valid = InputSplitter_io_Out_data_field1_0_valid; // @[extracted_function_reduction.scala 603:26]
  assign Loop_5_io_InLiveIn_11_bits_taskID = InputSplitter_io_Out_data_field1_0_bits_taskID; // @[extracted_function_reduction.scala 603:26]
  assign Loop_5_io_InLiveIn_11_bits_data = InputSplitter_io_Out_data_field1_0_bits_data; // @[extracted_function_reduction.scala 603:26]
  assign Loop_5_io_InLiveIn_12_valid = binaryOp_add125_io_Out_0_valid; // @[extracted_function_reduction.scala 605:26]
  assign Loop_5_io_InLiveIn_12_bits_data = binaryOp_add125_io_Out_0_bits_data; // @[extracted_function_reduction.scala 605:26]
  assign Loop_5_io_InLiveIn_13_valid = binaryOp_add43_io_Out_0_valid; // @[extracted_function_reduction.scala 607:26]
  assign Loop_5_io_InLiveIn_13_bits_data = binaryOp_add43_io_Out_0_bits_data; // @[extracted_function_reduction.scala 607:26]
  assign Loop_5_io_InLiveIn_14_valid = binaryOp_add0_io_Out_0_valid; // @[extracted_function_reduction.scala 609:26]
  assign Loop_5_io_InLiveIn_14_bits_data = binaryOp_add0_io_Out_0_bits_data; // @[extracted_function_reduction.scala 609:26]
  assign Loop_5_io_OutLiveIn_field14_0_ready = icmp_exitcond14817_io_RightIO_ready; // @[extracted_function_reduction.scala 669:33]
  assign Loop_5_io_OutLiveIn_field13_0_ready = Loop_4_io_InLiveIn_9_ready; // @[extracted_function_reduction.scala 575:25]
  assign Loop_5_io_OutLiveIn_field12_0_ready = Loop_4_io_InLiveIn_5_ready; // @[extracted_function_reduction.scala 567:25]
  assign Loop_5_io_OutLiveIn_field11_0_ready = Loop_4_io_InLiveIn_4_ready; // @[extracted_function_reduction.scala 565:25]
  assign Loop_5_io_OutLiveIn_field10_0_ready = Loop_4_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 559:25]
  assign Loop_5_io_OutLiveIn_field9_0_ready = Loop_4_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 561:25]
  assign Loop_5_io_OutLiveIn_field8_0_ready = Loop_4_io_InLiveIn_3_ready; // @[extracted_function_reduction.scala 563:25]
  assign Loop_5_io_OutLiveIn_field7_0_ready = Loop_4_io_InLiveIn_6_ready; // @[extracted_function_reduction.scala 569:25]
  assign Loop_5_io_OutLiveIn_field6_0_ready = Loop_4_io_InLiveIn_7_ready; // @[extracted_function_reduction.scala 571:25]
  assign Loop_5_io_OutLiveIn_field5_0_ready = Loop_4_io_InLiveIn_11_ready; // @[extracted_function_reduction.scala 579:26]
  assign Loop_5_io_OutLiveIn_field4_0_ready = Loop_4_io_InLiveIn_8_ready; // @[extracted_function_reduction.scala 573:25]
  assign Loop_5_io_OutLiveIn_field3_0_ready = Loop_4_io_InLiveIn_10_ready; // @[extracted_function_reduction.scala 577:26]
  assign Loop_5_io_OutLiveIn_field2_0_ready = br_13_io_CmpIO_ready; // @[extracted_function_reduction.scala 667:18]
  assign Loop_5_io_OutLiveIn_field1_0_ready = binaryOp_mul112_io_RightIO_ready; // @[extracted_function_reduction.scala 665:30]
  assign Loop_5_io_OutLiveIn_field0_0_ready = phi_pw_conv_reduction_s1_k_014310_io_InData_0_ready; // @[extracted_function_reduction.scala 661:50]
  assign Loop_5_io_OutLiveIn_field0_1_ready = binaryOp_sub11_io_RightIO_ready; // @[extracted_function_reduction.scala 663:29]
  assign Loop_5_io_activate_loop_start_ready = bb_for_body4_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 419:34]
  assign Loop_5_io_activate_loop_back_ready = bb_for_body4_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 421:34]
  assign Loop_5_io_loopBack_0_valid = br_18_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 497:25]
  assign Loop_5_io_loopBack_0_bits_taskID = br_18_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 497:25]
  assign Loop_5_io_loopBack_0_bits_control = br_18_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 497:25]
  assign Loop_5_io_loopFinish_0_valid = br_18_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 499:27]
  assign Loop_5_io_loopFinish_0_bits_control = br_18_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 499:27]
  assign Loop_5_io_CarryDepenIn_0_valid = binaryOp_inc6416_io_Out_0_valid; // @[extracted_function_reduction.scala 711:29]
  assign Loop_5_io_CarryDepenIn_0_bits_taskID = binaryOp_inc6416_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 711:29]
  assign Loop_5_io_CarryDepenIn_0_bits_data = binaryOp_inc6416_io_Out_0_bits_data; // @[extracted_function_reduction.scala 711:29]
  assign Loop_5_io_CarryDepenOut_field0_0_ready = phi_pw_conv_reduction_s1_k_014310_io_InData_1_ready; // @[extracted_function_reduction.scala 733:50]
  assign Loop_5_io_loopExit_0_ready = bb_for_cond_cleanup_loopexit2_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 417:51]
  assign bb_entry0_clock = clock;
  assign bb_entry0_reset = reset;
  assign bb_entry0_io_predicateIn_0_valid = InputSplitter_io_Out_enable_valid; // @[extracted_function_reduction.scala 391:31]
  assign bb_entry0_io_predicateIn_0_bits_taskID = InputSplitter_io_Out_enable_bits_taskID; // @[extracted_function_reduction.scala 391:31]
  assign bb_entry0_io_predicateIn_0_bits_control = InputSplitter_io_Out_enable_bits_control; // @[extracted_function_reduction.scala 391:31]
  assign bb_entry0_io_Out_0_ready = binaryOp_add0_io_enable_ready; // @[extracted_function_reduction.scala 741:27]
  assign bb_entry0_io_Out_1_ready = icmp_cmp1421_io_enable_ready; // @[extracted_function_reduction.scala 744:26]
  assign bb_entry0_io_Out_2_ready = br_2_io_enable_ready; // @[extracted_function_reduction.scala 747:18]
  assign bb_for_body_lr_ph1_clock = clock;
  assign bb_for_body_lr_ph1_reset = reset;
  assign bb_for_body_lr_ph1_io_predicateIn_0_valid = br_2_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 393:40]
  assign bb_for_body_lr_ph1_io_predicateIn_0_bits_taskID = br_2_io_TrueOutput_0_bits_taskID; // @[extracted_function_reduction.scala 393:40]
  assign bb_for_body_lr_ph1_io_predicateIn_0_bits_control = br_2_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 393:40]
  assign bb_for_body_lr_ph1_io_Out_0_ready = binaryOp_add43_io_enable_ready; // @[extracted_function_reduction.scala 750:28]
  assign bb_for_body_lr_ph1_io_Out_1_ready = icmp_cmp51394_io_enable_ready; // @[extracted_function_reduction.scala 753:27]
  assign bb_for_body_lr_ph1_io_Out_2_ready = binaryOp_add125_io_enable_ready; // @[extracted_function_reduction.scala 756:29]
  assign bb_for_body_lr_ph1_io_Out_3_ready = icmp_cmp131376_io_enable_ready; // @[extracted_function_reduction.scala 759:28]
  assign bb_for_body_lr_ph1_io_Out_4_ready = br_7_io_enable_ready; // @[extracted_function_reduction.scala 762:18]
  assign bb_for_cond_cleanup_loopexit2_clock = clock;
  assign bb_for_cond_cleanup_loopexit2_reset = reset;
  assign bb_for_cond_cleanup_loopexit2_io_predicateIn_0_valid = Loop_5_io_loopExit_0_valid; // @[extracted_function_reduction.scala 417:51]
  assign bb_for_cond_cleanup_loopexit2_io_predicateIn_0_bits_taskID = Loop_5_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 417:51]
  assign bb_for_cond_cleanup_loopexit2_io_predicateIn_0_bits_control = Loop_5_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 417:51]
  assign bb_for_cond_cleanup_loopexit2_io_Out_0_ready = br_8_io_enable_ready; // @[extracted_function_reduction.scala 765:18]
  assign bb_for_cond_cleanup3_clock = clock;
  assign bb_for_cond_cleanup3_reset = reset;
  assign bb_for_cond_cleanup3_io_predicateIn_0_valid = br_8_io_Out_0_valid; // @[extracted_function_reduction.scala 397:42]
  assign bb_for_cond_cleanup3_io_predicateIn_0_bits_taskID = br_8_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 397:42]
  assign bb_for_cond_cleanup3_io_predicateIn_0_bits_control = br_8_io_Out_0_bits_control; // @[extracted_function_reduction.scala 397:42]
  assign bb_for_cond_cleanup3_io_predicateIn_1_valid = br_2_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 395:42]
  assign bb_for_cond_cleanup3_io_predicateIn_1_bits_taskID = br_2_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 395:42]
  assign bb_for_cond_cleanup3_io_predicateIn_1_bits_control = br_2_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 395:42]
  assign bb_for_cond_cleanup3_io_Out_0_ready = ret_9_io_In_enable_ready; // @[extracted_function_reduction.scala 768:22]
  assign bb_for_body4_clock = clock;
  assign bb_for_body4_reset = reset;
  assign bb_for_body4_io_MaskBB_0_ready = phi_pw_conv_reduction_s1_k_014310_io_Mask_ready; // @[extracted_function_reduction.scala 988:45]
  assign bb_for_body4_io_Out_0_ready = phi_pw_conv_reduction_s1_k_014310_io_enable_ready; // @[extracted_function_reduction.scala 771:47]
  assign bb_for_body4_io_Out_1_ready = binaryOp_sub11_io_enable_ready; // @[extracted_function_reduction.scala 774:28]
  assign bb_for_body4_io_Out_2_ready = binaryOp_mul112_io_enable_ready; // @[extracted_function_reduction.scala 777:29]
  assign bb_for_body4_io_Out_3_ready = br_13_io_enable_ready; // @[extracted_function_reduction.scala 780:19]
  assign bb_for_body4_io_predicateIn_0_valid = Loop_5_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 421:34]
  assign bb_for_body4_io_predicateIn_0_bits_taskID = Loop_5_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 421:34]
  assign bb_for_body4_io_predicateIn_0_bits_control = Loop_5_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 421:34]
  assign bb_for_body4_io_predicateIn_1_valid = Loop_5_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 419:34]
  assign bb_for_body4_io_predicateIn_1_bits_taskID = Loop_5_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 419:34]
  assign bb_for_body4_io_predicateIn_1_bits_control = Loop_5_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 419:34]
  assign bb_for_body7_preheader5_clock = clock;
  assign bb_for_body7_preheader5_reset = reset;
  assign bb_for_body7_preheader5_io_predicateIn_0_valid = br_13_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 399:45]
  assign bb_for_body7_preheader5_io_predicateIn_0_bits_taskID = br_13_io_TrueOutput_0_bits_taskID; // @[extracted_function_reduction.scala 399:45]
  assign bb_for_body7_preheader5_io_predicateIn_0_bits_control = br_13_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 399:45]
  assign bb_for_body7_preheader5_io_Out_0_ready = br_14_io_enable_ready; // @[extracted_function_reduction.scala 783:19]
  assign bb_for_cond_cleanup6_loopexit6_clock = clock;
  assign bb_for_cond_cleanup6_loopexit6_reset = reset;
  assign bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_valid = Loop_4_io_loopExit_0_valid; // @[extracted_function_reduction.scala 423:52]
  assign bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_bits_taskID = Loop_4_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 423:52]
  assign bb_for_cond_cleanup6_loopexit6_io_predicateIn_0_bits_control = Loop_4_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 423:52]
  assign bb_for_cond_cleanup6_loopexit6_io_Out_0_ready = br_15_io_enable_ready; // @[extracted_function_reduction.scala 786:19]
  assign bb_for_cond_cleanup67_clock = clock;
  assign bb_for_cond_cleanup67_reset = reset;
  assign bb_for_cond_cleanup67_io_predicateIn_0_valid = br_15_io_Out_0_valid; // @[extracted_function_reduction.scala 403:43]
  assign bb_for_cond_cleanup67_io_predicateIn_0_bits_taskID = br_15_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 403:43]
  assign bb_for_cond_cleanup67_io_predicateIn_0_bits_control = br_15_io_Out_0_bits_control; // @[extracted_function_reduction.scala 403:43]
  assign bb_for_cond_cleanup67_io_predicateIn_1_valid = br_13_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 401:43]
  assign bb_for_cond_cleanup67_io_predicateIn_1_bits_taskID = br_13_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 401:43]
  assign bb_for_cond_cleanup67_io_predicateIn_1_bits_control = br_13_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 401:43]
  assign bb_for_cond_cleanup67_io_Out_0_ready = const0_io_enable_ready; // @[extracted_function_reduction.scala 789:20]
  assign bb_for_cond_cleanup67_io_Out_1_ready = binaryOp_inc6416_io_enable_ready; // @[extracted_function_reduction.scala 791:30]
  assign bb_for_cond_cleanup67_io_Out_2_ready = icmp_exitcond14817_io_enable_ready; // @[extracted_function_reduction.scala 794:32]
  assign bb_for_cond_cleanup67_io_Out_3_ready = br_18_io_enable_ready; // @[extracted_function_reduction.scala 797:19]
  assign bb_for_body78_clock = clock;
  assign bb_for_body78_reset = reset;
  assign bb_for_body78_io_MaskBB_0_ready = phi_pw_conv_reduction_s1_y_014019_io_Mask_ready; // @[extracted_function_reduction.scala 990:45]
  assign bb_for_body78_io_Out_0_ready = phi_pw_conv_reduction_s1_y_014019_io_enable_ready; // @[extracted_function_reduction.scala 800:47]
  assign bb_for_body78_io_Out_1_ready = br_20_io_enable_ready; // @[extracted_function_reduction.scala 803:19]
  assign bb_for_body78_io_predicateIn_0_valid = Loop_4_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 427:35]
  assign bb_for_body78_io_predicateIn_0_bits_taskID = Loop_4_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 427:35]
  assign bb_for_body78_io_predicateIn_0_bits_control = Loop_4_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 427:35]
  assign bb_for_body78_io_predicateIn_1_valid = Loop_4_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 425:35]
  assign bb_for_body78_io_predicateIn_1_bits_taskID = Loop_4_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 425:35]
  assign bb_for_body78_io_predicateIn_1_bits_control = Loop_4_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 425:35]
  assign bb_for_body15_lr_ph9_clock = clock;
  assign bb_for_body15_lr_ph9_reset = reset;
  assign bb_for_body15_lr_ph9_io_predicateIn_0_valid = br_20_io_TrueOutput_0_valid; // @[extracted_function_reduction.scala 405:42]
  assign bb_for_body15_lr_ph9_io_predicateIn_0_bits_taskID = br_20_io_TrueOutput_0_bits_taskID; // @[extracted_function_reduction.scala 405:42]
  assign bb_for_body15_lr_ph9_io_predicateIn_0_bits_control = br_20_io_TrueOutput_0_bits_control; // @[extracted_function_reduction.scala 405:42]
  assign bb_for_body15_lr_ph9_io_Out_0_ready = binaryOp_sub821_io_enable_ready; // @[extracted_function_reduction.scala 806:29]
  assign bb_for_body15_lr_ph9_io_Out_1_ready = binaryOp_reass_add22_io_enable_ready; // @[extracted_function_reduction.scala 809:34]
  assign bb_for_body15_lr_ph9_io_Out_2_ready = binaryOp_reass_mul23_io_enable_ready; // @[extracted_function_reduction.scala 812:34]
  assign bb_for_body15_lr_ph9_io_Out_3_ready = br_24_io_enable_ready; // @[extracted_function_reduction.scala 815:19]
  assign bb_for_cond_cleanup14_loopexit10_clock = clock;
  assign bb_for_cond_cleanup14_loopexit10_reset = reset;
  assign bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_valid = Loop_3_io_loopExit_0_valid; // @[extracted_function_reduction.scala 429:54]
  assign bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_bits_taskID = Loop_3_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 429:54]
  assign bb_for_cond_cleanup14_loopexit10_io_predicateIn_0_bits_control = Loop_3_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 429:54]
  assign bb_for_cond_cleanup14_loopexit10_io_Out_0_ready = br_25_io_enable_ready; // @[extracted_function_reduction.scala 818:19]
  assign bb_for_cond_cleanup1411_clock = clock;
  assign bb_for_cond_cleanup1411_reset = reset;
  assign bb_for_cond_cleanup1411_io_predicateIn_0_valid = br_25_io_Out_0_valid; // @[extracted_function_reduction.scala 409:45]
  assign bb_for_cond_cleanup1411_io_predicateIn_0_bits_taskID = br_25_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 409:45]
  assign bb_for_cond_cleanup1411_io_predicateIn_0_bits_control = br_25_io_Out_0_bits_control; // @[extracted_function_reduction.scala 409:45]
  assign bb_for_cond_cleanup1411_io_predicateIn_1_valid = br_20_io_FalseOutput_0_valid; // @[extracted_function_reduction.scala 407:45]
  assign bb_for_cond_cleanup1411_io_predicateIn_1_bits_taskID = br_20_io_FalseOutput_0_bits_taskID; // @[extracted_function_reduction.scala 407:45]
  assign bb_for_cond_cleanup1411_io_predicateIn_1_bits_control = br_20_io_FalseOutput_0_bits_control; // @[extracted_function_reduction.scala 407:45]
  assign bb_for_cond_cleanup1411_io_Out_0_ready = const1_io_enable_ready; // @[extracted_function_reduction.scala 821:20]
  assign bb_for_cond_cleanup1411_io_Out_1_ready = binaryOp_inc6126_io_enable_ready; // @[extracted_function_reduction.scala 823:30]
  assign bb_for_cond_cleanup1411_io_Out_2_ready = icmp_exitcond14727_io_enable_ready; // @[extracted_function_reduction.scala 826:32]
  assign bb_for_cond_cleanup1411_io_Out_3_ready = br_28_io_enable_ready; // @[extracted_function_reduction.scala 829:19]
  assign bb_for_body1512_clock = clock;
  assign bb_for_body1512_reset = reset;
  assign bb_for_body1512_io_MaskBB_0_ready = phi_pw_conv_reduction_s1_x_013829_io_Mask_ready; // @[extracted_function_reduction.scala 992:45]
  assign bb_for_body1512_io_Out_0_ready = phi_pw_conv_reduction_s1_x_013829_io_enable_ready; // @[extracted_function_reduction.scala 832:47]
  assign bb_for_body1512_io_Out_1_ready = binaryOp_sub1630_io_enable_ready; // @[extracted_function_reduction.scala 835:30]
  assign bb_for_body1512_io_Out_2_ready = binaryOp_add1031_io_enable_ready; // @[extracted_function_reduction.scala 838:30]
  assign bb_for_body1512_io_Out_3_ready = binaryOp_add1732_io_enable_ready; // @[extracted_function_reduction.scala 841:30]
  assign bb_for_body1512_io_Out_4_ready = Gep_arrayidx5033_io_enable_ready; // @[extracted_function_reduction.scala 844:30]
  assign bb_for_body1512_io_Out_5_ready = br_34_io_enable_ready; // @[extracted_function_reduction.scala 847:19]
  assign bb_for_body1512_io_predicateIn_0_valid = Loop_3_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 433:37]
  assign bb_for_body1512_io_predicateIn_0_bits_taskID = Loop_3_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 433:37]
  assign bb_for_body1512_io_predicateIn_0_bits_control = Loop_3_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 433:37]
  assign bb_for_body1512_io_predicateIn_1_valid = Loop_3_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 431:37]
  assign bb_for_body1512_io_predicateIn_1_bits_taskID = Loop_3_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 431:37]
  assign bb_for_body1512_io_predicateIn_1_bits_control = Loop_3_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 431:37]
  assign bb_for_cond_cleanup2013_clock = clock;
  assign bb_for_cond_cleanup2013_reset = reset;
  assign bb_for_cond_cleanup2013_io_predicateIn_0_valid = Loop_2_io_loopExit_0_valid; // @[extracted_function_reduction.scala 435:45]
  assign bb_for_cond_cleanup2013_io_predicateIn_0_bits_taskID = Loop_2_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 435:45]
  assign bb_for_cond_cleanup2013_io_predicateIn_0_bits_control = Loop_2_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 435:45]
  assign bb_for_cond_cleanup2013_io_Out_0_ready = const2_io_enable_ready; // @[extracted_function_reduction.scala 850:20]
  assign bb_for_cond_cleanup2013_io_Out_1_ready = binaryOp_inc5835_io_enable_ready; // @[extracted_function_reduction.scala 852:30]
  assign bb_for_cond_cleanup2013_io_Out_2_ready = icmp_exitcond14636_io_enable_ready; // @[extracted_function_reduction.scala 855:32]
  assign bb_for_cond_cleanup2013_io_Out_3_ready = br_37_io_enable_ready; // @[extracted_function_reduction.scala 858:19]
  assign bb_for_body2114_clock = clock;
  assign bb_for_body2114_reset = reset;
  assign bb_for_body2114_io_MaskBB_0_ready = phi_pw_conv_reduction_s1_r_pw__x_013638_io_Mask_ready; // @[extracted_function_reduction.scala 994:51]
  assign bb_for_body2114_io_Out_0_ready = const3_io_enable_ready; // @[extracted_function_reduction.scala 861:20]
  assign bb_for_body2114_io_Out_1_ready = phi_pw_conv_reduction_s1_r_pw__x_013638_io_enable_ready; // @[extracted_function_reduction.scala 863:53]
  assign bb_for_body2114_io_Out_2_ready = binaryOp_mul2239_io_enable_ready; // @[extracted_function_reduction.scala 866:30]
  assign bb_for_body2114_io_Out_3_ready = binaryOp_add2340_io_enable_ready; // @[extracted_function_reduction.scala 869:30]
  assign bb_for_body2114_io_Out_4_ready = br_41_io_enable_ready; // @[extracted_function_reduction.scala 872:19]
  assign bb_for_body2114_io_predicateIn_0_valid = Loop_2_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 439:37]
  assign bb_for_body2114_io_predicateIn_0_bits_taskID = Loop_2_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 439:37]
  assign bb_for_body2114_io_predicateIn_0_bits_control = Loop_2_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 439:37]
  assign bb_for_body2114_io_predicateIn_1_valid = Loop_2_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 437:37]
  assign bb_for_body2114_io_predicateIn_1_bits_taskID = Loop_2_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 437:37]
  assign bb_for_body2114_io_predicateIn_1_bits_control = Loop_2_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 437:37]
  assign bb_for_cond_cleanup2615_clock = clock;
  assign bb_for_cond_cleanup2615_reset = reset;
  assign bb_for_cond_cleanup2615_io_Out_0_ready = const4_io_enable_ready; // @[extracted_function_reduction.scala 875:20]
  assign bb_for_cond_cleanup2615_io_Out_1_ready = const5_io_enable_ready; // @[extracted_function_reduction.scala 877:20]
  assign bb_for_cond_cleanup2615_io_Out_2_ready = const6_io_enable_ready; // @[extracted_function_reduction.scala 879:20]
  assign bb_for_cond_cleanup2615_io_Out_3_ready = phiadd38_lcssa_lcssa42_io_enable_ready; // @[extracted_function_reduction.scala 881:36]
  assign bb_for_cond_cleanup2615_io_Out_4_ready = binaryOp_mul4443_io_enable_ready; // @[extracted_function_reduction.scala 884:30]
  assign bb_for_cond_cleanup2615_io_Out_5_ready = sextconv4744_io_enable_ready; // @[extracted_function_reduction.scala 887:26]
  assign bb_for_cond_cleanup2615_io_Out_6_ready = ld_45_io_enable_ready; // @[extracted_function_reduction.scala 890:19]
  assign bb_for_cond_cleanup2615_io_Out_7_ready = binaryOp_add5246_io_enable_ready; // @[extracted_function_reduction.scala 893:30]
  assign bb_for_cond_cleanup2615_io_Out_8_ready = st_47_io_enable_ready; // @[extracted_function_reduction.scala 896:19]
  assign bb_for_cond_cleanup2615_io_Out_9_ready = binaryOp_inc5548_io_enable_ready; // @[extracted_function_reduction.scala 899:30]
  assign bb_for_cond_cleanup2615_io_Out_10_ready = icmp_exitcond14549_io_enable_ready; // @[extracted_function_reduction.scala 902:32]
  assign bb_for_cond_cleanup2615_io_Out_11_ready = br_50_io_enable_ready; // @[extracted_function_reduction.scala 905:19]
  assign bb_for_cond_cleanup2615_io_predicateIn_0_valid = Loop_1_io_loopExit_0_valid; // @[extracted_function_reduction.scala 441:45]
  assign bb_for_cond_cleanup2615_io_predicateIn_0_bits_taskID = Loop_1_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 441:45]
  assign bb_for_cond_cleanup2615_io_predicateIn_0_bits_control = Loop_1_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 441:45]
  assign bb_for_body2716_clock = clock;
  assign bb_for_body2716_reset = reset;
  assign bb_for_body2716_io_MaskBB_0_ready = phi_dw_conv_013551_io_Mask_ready; // @[extracted_function_reduction.scala 998:30]
  assign bb_for_body2716_io_MaskBB_1_ready = phi_dw_conv_s1_r_dw__y_013452_io_Mask_ready; // @[extracted_function_reduction.scala 1000:41]
  assign bb_for_body2716_io_Out_0_ready = const7_io_enable_ready; // @[extracted_function_reduction.scala 908:20]
  assign bb_for_body2716_io_Out_1_ready = const8_io_enable_ready; // @[extracted_function_reduction.scala 910:20]
  assign bb_for_body2716_io_Out_2_ready = phi_dw_conv_013551_io_enable_ready; // @[extracted_function_reduction.scala 912:32]
  assign bb_for_body2716_io_Out_3_ready = phi_dw_conv_s1_r_dw__y_013452_io_enable_ready; // @[extracted_function_reduction.scala 915:43]
  assign bb_for_body2716_io_Out_4_ready = binaryOp_add2853_io_enable_ready; // @[extracted_function_reduction.scala 918:30]
  assign bb_for_body2716_io_Out_5_ready = binaryOp_mul2954_io_enable_ready; // @[extracted_function_reduction.scala 921:30]
  assign bb_for_body2716_io_Out_6_ready = binaryOp_add3055_io_enable_ready; // @[extracted_function_reduction.scala 924:30]
  assign bb_for_body2716_io_Out_7_ready = br_56_io_enable_ready; // @[extracted_function_reduction.scala 927:19]
  assign bb_for_body2716_io_predicateIn_0_valid = Loop_1_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 445:37]
  assign bb_for_body2716_io_predicateIn_0_bits_taskID = Loop_1_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 445:37]
  assign bb_for_body2716_io_predicateIn_0_bits_control = Loop_1_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 445:37]
  assign bb_for_body2716_io_predicateIn_1_valid = Loop_1_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 443:37]
  assign bb_for_body2716_io_predicateIn_1_bits_taskID = Loop_1_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 443:37]
  assign bb_for_body2716_io_predicateIn_1_bits_control = Loop_1_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 443:37]
  assign bb_for_cond_cleanup3317_clock = clock;
  assign bb_for_cond_cleanup3317_reset = reset;
  assign bb_for_cond_cleanup3317_io_Out_0_ready = const9_io_enable_ready; // @[extracted_function_reduction.scala 930:20]
  assign bb_for_cond_cleanup3317_io_Out_1_ready = const10_io_enable_ready; // @[extracted_function_reduction.scala 932:21]
  assign bb_for_cond_cleanup3317_io_Out_2_ready = phiadd38_lcssa57_io_enable_ready; // @[extracted_function_reduction.scala 934:30]
  assign bb_for_cond_cleanup3317_io_Out_3_ready = binaryOp_inc4158_io_enable_ready; // @[extracted_function_reduction.scala 937:30]
  assign bb_for_cond_cleanup3317_io_Out_4_ready = icmp_exitcond14459_io_enable_ready; // @[extracted_function_reduction.scala 940:32]
  assign bb_for_cond_cleanup3317_io_Out_5_ready = br_60_io_enable_ready; // @[extracted_function_reduction.scala 943:19]
  assign bb_for_cond_cleanup3317_io_predicateIn_0_valid = Loop_0_io_loopExit_0_valid; // @[extracted_function_reduction.scala 447:45]
  assign bb_for_cond_cleanup3317_io_predicateIn_0_bits_taskID = Loop_0_io_loopExit_0_bits_taskID; // @[extracted_function_reduction.scala 447:45]
  assign bb_for_cond_cleanup3317_io_predicateIn_0_bits_control = Loop_0_io_loopExit_0_bits_control; // @[extracted_function_reduction.scala 447:45]
  assign bb_for_body3418_clock = clock;
  assign bb_for_body3418_reset = reset;
  assign bb_for_body3418_io_MaskBB_0_ready = phi_dw_conv_113361_io_Mask_ready; // @[extracted_function_reduction.scala 1004:30]
  assign bb_for_body3418_io_MaskBB_1_ready = phi_dw_conv_s1_r_dw__x_013262_io_Mask_ready; // @[extracted_function_reduction.scala 1006:41]
  assign bb_for_body3418_io_Out_0_ready = const11_io_enable_ready; // @[extracted_function_reduction.scala 946:21]
  assign bb_for_body3418_io_Out_1_ready = const12_io_enable_ready; // @[extracted_function_reduction.scala 948:21]
  assign bb_for_body3418_io_Out_2_ready = const13_io_enable_ready; // @[extracted_function_reduction.scala 950:21]
  assign bb_for_body3418_io_Out_3_ready = phi_dw_conv_113361_io_enable_ready; // @[extracted_function_reduction.scala 952:32]
  assign bb_for_body3418_io_Out_4_ready = phi_dw_conv_s1_r_dw__x_013262_io_enable_ready; // @[extracted_function_reduction.scala 955:43]
  assign bb_for_body3418_io_Out_5_ready = binaryOp_add3563_io_enable_ready; // @[extracted_function_reduction.scala 958:30]
  assign bb_for_body3418_io_Out_6_ready = Gep_arrayidx64_io_enable_ready; // @[extracted_function_reduction.scala 961:28]
  assign bb_for_body3418_io_Out_7_ready = ld_65_io_enable_ready; // @[extracted_function_reduction.scala 964:19]
  assign bb_for_body3418_io_Out_8_ready = sextconv3766_io_enable_ready; // @[extracted_function_reduction.scala 967:26]
  assign bb_for_body3418_io_Out_9_ready = binaryOp_add3867_io_enable_ready; // @[extracted_function_reduction.scala 970:30]
  assign bb_for_body3418_io_Out_10_ready = binaryOp_inc68_io_enable_ready; // @[extracted_function_reduction.scala 973:28]
  assign bb_for_body3418_io_Out_11_ready = icmp_exitcond69_io_enable_ready; // @[extracted_function_reduction.scala 976:29]
  assign bb_for_body3418_io_Out_12_ready = br_70_io_enable_ready; // @[extracted_function_reduction.scala 979:19]
  assign bb_for_body3418_io_predicateIn_0_valid = Loop_0_io_activate_loop_back_valid; // @[extracted_function_reduction.scala 451:37]
  assign bb_for_body3418_io_predicateIn_0_bits_taskID = Loop_0_io_activate_loop_back_bits_taskID; // @[extracted_function_reduction.scala 451:37]
  assign bb_for_body3418_io_predicateIn_0_bits_control = Loop_0_io_activate_loop_back_bits_control; // @[extracted_function_reduction.scala 451:37]
  assign bb_for_body3418_io_predicateIn_1_valid = Loop_0_io_activate_loop_start_valid; // @[extracted_function_reduction.scala 449:37]
  assign bb_for_body3418_io_predicateIn_1_bits_taskID = Loop_0_io_activate_loop_start_bits_taskID; // @[extracted_function_reduction.scala 449:37]
  assign bb_for_body3418_io_predicateIn_1_bits_control = Loop_0_io_activate_loop_start_bits_control; // @[extracted_function_reduction.scala 449:37]
  assign binaryOp_add0_clock = clock;
  assign binaryOp_add0_reset = reset;
  assign binaryOp_add0_io_enable_valid = bb_entry0_io_Out_0_valid; // @[extracted_function_reduction.scala 741:27]
  assign binaryOp_add0_io_enable_bits_taskID = bb_entry0_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 741:27]
  assign binaryOp_add0_io_enable_bits_control = bb_entry0_io_Out_0_bits_control; // @[extracted_function_reduction.scala 741:27]
  assign binaryOp_add0_io_Out_0_ready = Loop_5_io_InLiveIn_14_ready; // @[extracted_function_reduction.scala 609:26]
  assign binaryOp_add0_io_Out_1_ready = icmp_cmp1421_io_LeftIO_ready; // @[extracted_function_reduction.scala 1072:26]
  assign binaryOp_add0_io_LeftIO_valid = InputSplitter_io_Out_data_field9_0_valid; // @[extracted_function_reduction.scala 1182:27]
  assign binaryOp_add0_io_LeftIO_bits_data = InputSplitter_io_Out_data_field9_0_bits_data; // @[extracted_function_reduction.scala 1182:27]
  assign binaryOp_add0_io_RightIO_valid = InputSplitter_io_Out_data_field8_1_valid; // @[extracted_function_reduction.scala 1178:28]
  assign binaryOp_add0_io_RightIO_bits_data = InputSplitter_io_Out_data_field8_1_bits_data; // @[extracted_function_reduction.scala 1178:28]
  assign icmp_cmp1421_clock = clock;
  assign icmp_cmp1421_reset = reset;
  assign icmp_cmp1421_io_enable_valid = bb_entry0_io_Out_1_valid; // @[extracted_function_reduction.scala 744:26]
  assign icmp_cmp1421_io_enable_bits_taskID = bb_entry0_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 744:26]
  assign icmp_cmp1421_io_enable_bits_control = bb_entry0_io_Out_1_bits_control; // @[extracted_function_reduction.scala 744:26]
  assign icmp_cmp1421_io_Out_0_ready = br_2_io_CmpIO_ready; // @[extracted_function_reduction.scala 1074:17]
  assign icmp_cmp1421_io_LeftIO_valid = binaryOp_add0_io_Out_1_valid; // @[extracted_function_reduction.scala 1072:26]
  assign icmp_cmp1421_io_LeftIO_bits_data = binaryOp_add0_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1072:26]
  assign icmp_cmp1421_io_RightIO_valid = InputSplitter_io_Out_data_field8_2_valid; // @[extracted_function_reduction.scala 1180:27]
  assign icmp_cmp1421_io_RightIO_bits_data = InputSplitter_io_Out_data_field8_2_bits_data; // @[extracted_function_reduction.scala 1180:27]
  assign br_2_clock = clock;
  assign br_2_reset = reset;
  assign br_2_io_enable_valid = bb_entry0_io_Out_2_valid; // @[extracted_function_reduction.scala 747:18]
  assign br_2_io_enable_bits_taskID = bb_entry0_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 747:18]
  assign br_2_io_enable_bits_control = bb_entry0_io_Out_2_bits_control; // @[extracted_function_reduction.scala 747:18]
  assign br_2_io_CmpIO_valid = icmp_cmp1421_io_Out_0_valid; // @[extracted_function_reduction.scala 1074:17]
  assign br_2_io_CmpIO_bits_taskID = icmp_cmp1421_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 1074:17]
  assign br_2_io_CmpIO_bits_data = icmp_cmp1421_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1074:17]
  assign br_2_io_TrueOutput_0_ready = bb_for_body_lr_ph1_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 393:40]
  assign br_2_io_FalseOutput_0_ready = bb_for_cond_cleanup3_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 395:42]
  assign binaryOp_add43_clock = clock;
  assign binaryOp_add43_reset = reset;
  assign binaryOp_add43_io_enable_valid = bb_for_body_lr_ph1_io_Out_0_valid; // @[extracted_function_reduction.scala 750:28]
  assign binaryOp_add43_io_enable_bits_taskID = bb_for_body_lr_ph1_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 750:28]
  assign binaryOp_add43_io_enable_bits_control = bb_for_body_lr_ph1_io_Out_0_bits_control; // @[extracted_function_reduction.scala 750:28]
  assign binaryOp_add43_io_Out_0_ready = Loop_5_io_InLiveIn_13_ready; // @[extracted_function_reduction.scala 607:26]
  assign binaryOp_add43_io_Out_1_ready = icmp_cmp51394_io_LeftIO_ready; // @[extracted_function_reduction.scala 1076:27]
  assign binaryOp_add43_io_LeftIO_valid = InputSplitter_io_Out_data_field7_1_valid; // @[extracted_function_reduction.scala 1176:28]
  assign binaryOp_add43_io_LeftIO_bits_data = InputSplitter_io_Out_data_field7_1_bits_data; // @[extracted_function_reduction.scala 1176:28]
  assign binaryOp_add43_io_RightIO_valid = InputSplitter_io_Out_data_field6_1_valid; // @[extracted_function_reduction.scala 1172:29]
  assign binaryOp_add43_io_RightIO_bits_data = InputSplitter_io_Out_data_field6_1_bits_data; // @[extracted_function_reduction.scala 1172:29]
  assign icmp_cmp51394_clock = clock;
  assign icmp_cmp51394_reset = reset;
  assign icmp_cmp51394_io_enable_valid = bb_for_body_lr_ph1_io_Out_1_valid; // @[extracted_function_reduction.scala 753:27]
  assign icmp_cmp51394_io_enable_bits_taskID = bb_for_body_lr_ph1_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 753:27]
  assign icmp_cmp51394_io_enable_bits_control = bb_for_body_lr_ph1_io_Out_1_bits_control; // @[extracted_function_reduction.scala 753:27]
  assign icmp_cmp51394_io_Out_0_ready = Loop_5_io_InLiveIn_2_ready; // @[extracted_function_reduction.scala 585:25]
  assign icmp_cmp51394_io_LeftIO_valid = binaryOp_add43_io_Out_1_valid; // @[extracted_function_reduction.scala 1076:27]
  assign icmp_cmp51394_io_LeftIO_bits_data = binaryOp_add43_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1076:27]
  assign icmp_cmp51394_io_RightIO_valid = InputSplitter_io_Out_data_field6_2_valid; // @[extracted_function_reduction.scala 1174:28]
  assign icmp_cmp51394_io_RightIO_bits_data = InputSplitter_io_Out_data_field6_2_bits_data; // @[extracted_function_reduction.scala 1174:28]
  assign binaryOp_add125_clock = clock;
  assign binaryOp_add125_reset = reset;
  assign binaryOp_add125_io_enable_valid = bb_for_body_lr_ph1_io_Out_2_valid; // @[extracted_function_reduction.scala 756:29]
  assign binaryOp_add125_io_enable_bits_taskID = bb_for_body_lr_ph1_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 756:29]
  assign binaryOp_add125_io_enable_bits_control = bb_for_body_lr_ph1_io_Out_2_bits_control; // @[extracted_function_reduction.scala 756:29]
  assign binaryOp_add125_io_Out_0_ready = Loop_5_io_InLiveIn_12_ready; // @[extracted_function_reduction.scala 605:26]
  assign binaryOp_add125_io_Out_1_ready = icmp_cmp131376_io_LeftIO_ready; // @[extracted_function_reduction.scala 1078:28]
  assign binaryOp_add125_io_LeftIO_valid = InputSplitter_io_Out_data_field5_1_valid; // @[extracted_function_reduction.scala 1170:29]
  assign binaryOp_add125_io_LeftIO_bits_data = InputSplitter_io_Out_data_field5_1_bits_data; // @[extracted_function_reduction.scala 1170:29]
  assign binaryOp_add125_io_RightIO_valid = InputSplitter_io_Out_data_field4_1_valid; // @[extracted_function_reduction.scala 1166:30]
  assign binaryOp_add125_io_RightIO_bits_data = InputSplitter_io_Out_data_field4_1_bits_data; // @[extracted_function_reduction.scala 1166:30]
  assign icmp_cmp131376_clock = clock;
  assign icmp_cmp131376_reset = reset;
  assign icmp_cmp131376_io_enable_valid = bb_for_body_lr_ph1_io_Out_3_valid; // @[extracted_function_reduction.scala 759:28]
  assign icmp_cmp131376_io_enable_bits_taskID = bb_for_body_lr_ph1_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 759:28]
  assign icmp_cmp131376_io_enable_bits_control = bb_for_body_lr_ph1_io_Out_3_bits_control; // @[extracted_function_reduction.scala 759:28]
  assign icmp_cmp131376_io_Out_0_ready = Loop_5_io_InLiveIn_4_ready; // @[extracted_function_reduction.scala 589:25]
  assign icmp_cmp131376_io_LeftIO_valid = binaryOp_add125_io_Out_1_valid; // @[extracted_function_reduction.scala 1078:28]
  assign icmp_cmp131376_io_LeftIO_bits_data = binaryOp_add125_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1078:28]
  assign icmp_cmp131376_io_RightIO_valid = InputSplitter_io_Out_data_field4_2_valid; // @[extracted_function_reduction.scala 1168:29]
  assign icmp_cmp131376_io_RightIO_bits_data = InputSplitter_io_Out_data_field4_2_bits_data; // @[extracted_function_reduction.scala 1168:29]
  assign br_7_clock = clock;
  assign br_7_reset = reset;
  assign br_7_io_enable_valid = bb_for_body_lr_ph1_io_Out_4_valid; // @[extracted_function_reduction.scala 762:18]
  assign br_7_io_enable_bits_taskID = bb_for_body_lr_ph1_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 762:18]
  assign br_7_io_enable_bits_control = bb_for_body_lr_ph1_io_Out_4_bits_control; // @[extracted_function_reduction.scala 762:18]
  assign br_7_io_Out_0_ready = Loop_5_io_enable_ready; // @[extracted_function_reduction.scala 495:20]
  assign br_8_clock = clock;
  assign br_8_reset = reset;
  assign br_8_io_enable_valid = bb_for_cond_cleanup_loopexit2_io_Out_0_valid; // @[extracted_function_reduction.scala 765:18]
  assign br_8_io_enable_bits_taskID = bb_for_cond_cleanup_loopexit2_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 765:18]
  assign br_8_io_enable_bits_control = bb_for_cond_cleanup_loopexit2_io_Out_0_bits_control; // @[extracted_function_reduction.scala 765:18]
  assign br_8_io_Out_0_ready = bb_for_cond_cleanup3_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 397:42]
  assign ret_9_clock = clock;
  assign ret_9_reset = reset;
  assign ret_9_io_In_enable_valid = bb_for_cond_cleanup3_io_Out_0_valid; // @[extracted_function_reduction.scala 768:22]
  assign ret_9_io_In_enable_bits_taskID = bb_for_cond_cleanup3_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 768:22]
  assign ret_9_io_In_enable_bits_control = bb_for_cond_cleanup3_io_Out_0_bits_control; // @[extracted_function_reduction.scala 768:22]
  assign ret_9_io_Out_ready = io_out_ready; // @[extracted_function_reduction.scala 1192:10]
  assign phi_pw_conv_reduction_s1_k_014310_clock = clock;
  assign phi_pw_conv_reduction_s1_k_014310_reset = reset;
  assign phi_pw_conv_reduction_s1_k_014310_io_enable_valid = bb_for_body4_io_Out_0_valid; // @[extracted_function_reduction.scala 771:47]
  assign phi_pw_conv_reduction_s1_k_014310_io_enable_bits_control = bb_for_body4_io_Out_0_bits_control; // @[extracted_function_reduction.scala 771:47]
  assign phi_pw_conv_reduction_s1_k_014310_io_InData_0_valid = Loop_5_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 661:50]
  assign phi_pw_conv_reduction_s1_k_014310_io_InData_0_bits_taskID = Loop_5_io_OutLiveIn_field0_0_bits_taskID; // @[extracted_function_reduction.scala 661:50]
  assign phi_pw_conv_reduction_s1_k_014310_io_InData_0_bits_data = Loop_5_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 661:50]
  assign phi_pw_conv_reduction_s1_k_014310_io_InData_1_valid = Loop_5_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 733:50]
  assign phi_pw_conv_reduction_s1_k_014310_io_InData_1_bits_taskID = Loop_5_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 733:50]
  assign phi_pw_conv_reduction_s1_k_014310_io_InData_1_bits_data = Loop_5_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 733:50]
  assign phi_pw_conv_reduction_s1_k_014310_io_Mask_valid = bb_for_body4_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 988:45]
  assign phi_pw_conv_reduction_s1_k_014310_io_Mask_bits = bb_for_body4_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 988:45]
  assign phi_pw_conv_reduction_s1_k_014310_io_Out_0_ready = binaryOp_sub11_io_LeftIO_ready; // @[extracted_function_reduction.scala 1080:28]
  assign phi_pw_conv_reduction_s1_k_014310_io_Out_1_ready = binaryOp_inc6416_io_LeftIO_ready; // @[extracted_function_reduction.scala 1082:30]
  assign binaryOp_sub11_clock = clock;
  assign binaryOp_sub11_reset = reset;
  assign binaryOp_sub11_io_enable_valid = bb_for_body4_io_Out_1_valid; // @[extracted_function_reduction.scala 774:28]
  assign binaryOp_sub11_io_enable_bits_taskID = bb_for_body4_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 774:28]
  assign binaryOp_sub11_io_enable_bits_control = bb_for_body4_io_Out_1_bits_control; // @[extracted_function_reduction.scala 774:28]
  assign binaryOp_sub11_io_Out_0_ready = binaryOp_mul112_io_LeftIO_ready; // @[extracted_function_reduction.scala 1084:29]
  assign binaryOp_sub11_io_LeftIO_valid = phi_pw_conv_reduction_s1_k_014310_io_Out_0_valid; // @[extracted_function_reduction.scala 1080:28]
  assign binaryOp_sub11_io_LeftIO_bits_data = phi_pw_conv_reduction_s1_k_014310_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1080:28]
  assign binaryOp_sub11_io_RightIO_valid = Loop_5_io_OutLiveIn_field0_1_valid; // @[extracted_function_reduction.scala 663:29]
  assign binaryOp_sub11_io_RightIO_bits_data = Loop_5_io_OutLiveIn_field0_1_bits_data; // @[extracted_function_reduction.scala 663:29]
  assign binaryOp_mul112_clock = clock;
  assign binaryOp_mul112_reset = reset;
  assign binaryOp_mul112_io_enable_valid = bb_for_body4_io_Out_2_valid; // @[extracted_function_reduction.scala 777:29]
  assign binaryOp_mul112_io_enable_bits_taskID = bb_for_body4_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 777:29]
  assign binaryOp_mul112_io_enable_bits_control = bb_for_body4_io_Out_2_bits_control; // @[extracted_function_reduction.scala 777:29]
  assign binaryOp_mul112_io_Out_0_ready = Loop_4_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 557:25]
  assign binaryOp_mul112_io_LeftIO_valid = binaryOp_sub11_io_Out_0_valid; // @[extracted_function_reduction.scala 1084:29]
  assign binaryOp_mul112_io_LeftIO_bits_data = binaryOp_sub11_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1084:29]
  assign binaryOp_mul112_io_RightIO_valid = Loop_5_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 665:30]
  assign binaryOp_mul112_io_RightIO_bits_data = Loop_5_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 665:30]
  assign br_13_clock = clock;
  assign br_13_reset = reset;
  assign br_13_io_enable_valid = bb_for_body4_io_Out_3_valid; // @[extracted_function_reduction.scala 780:19]
  assign br_13_io_enable_bits_taskID = bb_for_body4_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 780:19]
  assign br_13_io_enable_bits_control = bb_for_body4_io_Out_3_bits_control; // @[extracted_function_reduction.scala 780:19]
  assign br_13_io_CmpIO_valid = Loop_5_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 667:18]
  assign br_13_io_CmpIO_bits_taskID = Loop_5_io_OutLiveIn_field2_0_bits_taskID; // @[extracted_function_reduction.scala 667:18]
  assign br_13_io_CmpIO_bits_data = Loop_5_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 667:18]
  assign br_13_io_TrueOutput_0_ready = bb_for_body7_preheader5_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 399:45]
  assign br_13_io_FalseOutput_0_ready = bb_for_cond_cleanup67_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 401:43]
  assign br_14_clock = clock;
  assign br_14_reset = reset;
  assign br_14_io_enable_valid = bb_for_body7_preheader5_io_Out_0_valid; // @[extracted_function_reduction.scala 783:19]
  assign br_14_io_enable_bits_taskID = bb_for_body7_preheader5_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 783:19]
  assign br_14_io_enable_bits_control = bb_for_body7_preheader5_io_Out_0_bits_control; // @[extracted_function_reduction.scala 783:19]
  assign br_14_io_Out_0_ready = Loop_4_io_enable_ready; // @[extracted_function_reduction.scala 489:20]
  assign br_15_clock = clock;
  assign br_15_reset = reset;
  assign br_15_io_enable_valid = bb_for_cond_cleanup6_loopexit6_io_Out_0_valid; // @[extracted_function_reduction.scala 786:19]
  assign br_15_io_enable_bits_taskID = bb_for_cond_cleanup6_loopexit6_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 786:19]
  assign br_15_io_enable_bits_control = bb_for_cond_cleanup6_loopexit6_io_Out_0_bits_control; // @[extracted_function_reduction.scala 786:19]
  assign br_15_io_Out_0_ready = bb_for_cond_cleanup67_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 403:43]
  assign binaryOp_inc6416_clock = clock;
  assign binaryOp_inc6416_reset = reset;
  assign binaryOp_inc6416_io_enable_valid = bb_for_cond_cleanup67_io_Out_1_valid; // @[extracted_function_reduction.scala 791:30]
  assign binaryOp_inc6416_io_enable_bits_taskID = bb_for_cond_cleanup67_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 791:30]
  assign binaryOp_inc6416_io_enable_bits_control = bb_for_cond_cleanup67_io_Out_1_bits_control; // @[extracted_function_reduction.scala 791:30]
  assign binaryOp_inc6416_io_Out_0_ready = Loop_5_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 711:29]
  assign binaryOp_inc6416_io_Out_1_ready = icmp_exitcond14817_io_LeftIO_ready; // @[extracted_function_reduction.scala 1086:32]
  assign binaryOp_inc6416_io_LeftIO_valid = phi_pw_conv_reduction_s1_k_014310_io_Out_1_valid; // @[extracted_function_reduction.scala 1082:30]
  assign binaryOp_inc6416_io_LeftIO_bits_data = phi_pw_conv_reduction_s1_k_014310_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1082:30]
  assign binaryOp_inc6416_io_RightIO_valid = const0_io_Out_valid; // @[extracted_function_reduction.scala 1044:31]
  assign icmp_exitcond14817_clock = clock;
  assign icmp_exitcond14817_reset = reset;
  assign icmp_exitcond14817_io_enable_valid = bb_for_cond_cleanup67_io_Out_2_valid; // @[extracted_function_reduction.scala 794:32]
  assign icmp_exitcond14817_io_enable_bits_taskID = bb_for_cond_cleanup67_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 794:32]
  assign icmp_exitcond14817_io_enable_bits_control = bb_for_cond_cleanup67_io_Out_2_bits_control; // @[extracted_function_reduction.scala 794:32]
  assign icmp_exitcond14817_io_Out_0_ready = br_18_io_CmpIO_ready; // @[extracted_function_reduction.scala 1088:18]
  assign icmp_exitcond14817_io_LeftIO_valid = binaryOp_inc6416_io_Out_1_valid; // @[extracted_function_reduction.scala 1086:32]
  assign icmp_exitcond14817_io_LeftIO_bits_data = binaryOp_inc6416_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1086:32]
  assign icmp_exitcond14817_io_RightIO_valid = Loop_5_io_OutLiveIn_field14_0_valid; // @[extracted_function_reduction.scala 669:33]
  assign icmp_exitcond14817_io_RightIO_bits_data = Loop_5_io_OutLiveIn_field14_0_bits_data; // @[extracted_function_reduction.scala 669:33]
  assign br_18_clock = clock;
  assign br_18_reset = reset;
  assign br_18_io_enable_valid = bb_for_cond_cleanup67_io_Out_3_valid; // @[extracted_function_reduction.scala 797:19]
  assign br_18_io_enable_bits_taskID = bb_for_cond_cleanup67_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 797:19]
  assign br_18_io_enable_bits_control = bb_for_cond_cleanup67_io_Out_3_bits_control; // @[extracted_function_reduction.scala 797:19]
  assign br_18_io_CmpIO_valid = icmp_exitcond14817_io_Out_0_valid; // @[extracted_function_reduction.scala 1088:18]
  assign br_18_io_CmpIO_bits_taskID = icmp_exitcond14817_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 1088:18]
  assign br_18_io_CmpIO_bits_data = icmp_exitcond14817_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1088:18]
  assign br_18_io_TrueOutput_0_ready = Loop_5_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 499:27]
  assign br_18_io_FalseOutput_0_ready = Loop_5_io_loopBack_0_ready; // @[extracted_function_reduction.scala 497:25]
  assign phi_pw_conv_reduction_s1_y_014019_clock = clock;
  assign phi_pw_conv_reduction_s1_y_014019_reset = reset;
  assign phi_pw_conv_reduction_s1_y_014019_io_enable_valid = bb_for_body78_io_Out_0_valid; // @[extracted_function_reduction.scala 800:47]
  assign phi_pw_conv_reduction_s1_y_014019_io_enable_bits_control = bb_for_body78_io_Out_0_bits_control; // @[extracted_function_reduction.scala 800:47]
  assign phi_pw_conv_reduction_s1_y_014019_io_InData_0_valid = Loop_4_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 731:50]
  assign phi_pw_conv_reduction_s1_y_014019_io_InData_0_bits_taskID = Loop_4_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 731:50]
  assign phi_pw_conv_reduction_s1_y_014019_io_InData_0_bits_data = Loop_4_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 731:50]
  assign phi_pw_conv_reduction_s1_y_014019_io_InData_1_valid = Loop_4_io_OutLiveIn_field10_0_valid; // @[extracted_function_reduction.scala 655:50]
  assign phi_pw_conv_reduction_s1_y_014019_io_InData_1_bits_taskID = Loop_4_io_OutLiveIn_field10_0_bits_taskID; // @[extracted_function_reduction.scala 655:50]
  assign phi_pw_conv_reduction_s1_y_014019_io_InData_1_bits_data = Loop_4_io_OutLiveIn_field10_0_bits_data; // @[extracted_function_reduction.scala 655:50]
  assign phi_pw_conv_reduction_s1_y_014019_io_Mask_valid = bb_for_body78_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 990:45]
  assign phi_pw_conv_reduction_s1_y_014019_io_Mask_bits = bb_for_body78_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 990:45]
  assign phi_pw_conv_reduction_s1_y_014019_io_Out_0_ready = Loop_3_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 541:25]
  assign phi_pw_conv_reduction_s1_y_014019_io_Out_1_ready = binaryOp_sub821_io_LeftIO_ready; // @[extracted_function_reduction.scala 1090:29]
  assign phi_pw_conv_reduction_s1_y_014019_io_Out_2_ready = binaryOp_inc6126_io_LeftIO_ready; // @[extracted_function_reduction.scala 1092:30]
  assign br_20_clock = clock;
  assign br_20_reset = reset;
  assign br_20_io_enable_valid = bb_for_body78_io_Out_1_valid; // @[extracted_function_reduction.scala 803:19]
  assign br_20_io_enable_bits_taskID = bb_for_body78_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 803:19]
  assign br_20_io_enable_bits_control = bb_for_body78_io_Out_1_bits_control; // @[extracted_function_reduction.scala 803:19]
  assign br_20_io_CmpIO_valid = Loop_4_io_OutLiveIn_field8_0_valid; // @[extracted_function_reduction.scala 651:18]
  assign br_20_io_CmpIO_bits_taskID = Loop_4_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_reduction.scala 651:18]
  assign br_20_io_CmpIO_bits_data = Loop_4_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_reduction.scala 651:18]
  assign br_20_io_TrueOutput_0_ready = bb_for_body15_lr_ph9_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 405:42]
  assign br_20_io_FalseOutput_0_ready = bb_for_cond_cleanup1411_io_predicateIn_1_ready; // @[extracted_function_reduction.scala 407:45]
  assign binaryOp_sub821_clock = clock;
  assign binaryOp_sub821_reset = reset;
  assign binaryOp_sub821_io_enable_valid = bb_for_body15_lr_ph9_io_Out_0_valid; // @[extracted_function_reduction.scala 806:29]
  assign binaryOp_sub821_io_enable_bits_taskID = bb_for_body15_lr_ph9_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 806:29]
  assign binaryOp_sub821_io_enable_bits_control = bb_for_body15_lr_ph9_io_Out_0_bits_control; // @[extracted_function_reduction.scala 806:29]
  assign binaryOp_sub821_io_Out_0_ready = binaryOp_reass_add22_io_LeftIO_ready; // @[extracted_function_reduction.scala 1094:34]
  assign binaryOp_sub821_io_LeftIO_valid = phi_pw_conv_reduction_s1_y_014019_io_Out_1_valid; // @[extracted_function_reduction.scala 1090:29]
  assign binaryOp_sub821_io_LeftIO_bits_data = phi_pw_conv_reduction_s1_y_014019_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1090:29]
  assign binaryOp_sub821_io_RightIO_valid = Loop_4_io_OutLiveIn_field10_1_valid; // @[extracted_function_reduction.scala 657:30]
  assign binaryOp_sub821_io_RightIO_bits_data = Loop_4_io_OutLiveIn_field10_1_bits_data; // @[extracted_function_reduction.scala 657:30]
  assign binaryOp_reass_add22_clock = clock;
  assign binaryOp_reass_add22_reset = reset;
  assign binaryOp_reass_add22_io_enable_valid = bb_for_body15_lr_ph9_io_Out_1_valid; // @[extracted_function_reduction.scala 809:34]
  assign binaryOp_reass_add22_io_enable_bits_taskID = bb_for_body15_lr_ph9_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 809:34]
  assign binaryOp_reass_add22_io_enable_bits_control = bb_for_body15_lr_ph9_io_Out_1_bits_control; // @[extracted_function_reduction.scala 809:34]
  assign binaryOp_reass_add22_io_Out_0_ready = binaryOp_reass_mul23_io_LeftIO_ready; // @[extracted_function_reduction.scala 1096:34]
  assign binaryOp_reass_add22_io_LeftIO_valid = binaryOp_sub821_io_Out_0_valid; // @[extracted_function_reduction.scala 1094:34]
  assign binaryOp_reass_add22_io_LeftIO_bits_data = binaryOp_sub821_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1094:34]
  assign binaryOp_reass_add22_io_RightIO_valid = Loop_4_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 649:35]
  assign binaryOp_reass_add22_io_RightIO_bits_data = Loop_4_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 649:35]
  assign binaryOp_reass_mul23_clock = clock;
  assign binaryOp_reass_mul23_reset = reset;
  assign binaryOp_reass_mul23_io_enable_valid = bb_for_body15_lr_ph9_io_Out_2_valid; // @[extracted_function_reduction.scala 812:34]
  assign binaryOp_reass_mul23_io_enable_bits_taskID = bb_for_body15_lr_ph9_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 812:34]
  assign binaryOp_reass_mul23_io_enable_bits_control = bb_for_body15_lr_ph9_io_Out_2_bits_control; // @[extracted_function_reduction.scala 812:34]
  assign binaryOp_reass_mul23_io_Out_0_ready = Loop_3_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 539:25]
  assign binaryOp_reass_mul23_io_LeftIO_valid = binaryOp_reass_add22_io_Out_0_valid; // @[extracted_function_reduction.scala 1096:34]
  assign binaryOp_reass_mul23_io_LeftIO_bits_data = binaryOp_reass_add22_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1096:34]
  assign binaryOp_reass_mul23_io_RightIO_valid = Loop_4_io_OutLiveIn_field11_0_valid; // @[extracted_function_reduction.scala 659:35]
  assign binaryOp_reass_mul23_io_RightIO_bits_data = Loop_4_io_OutLiveIn_field11_0_bits_data; // @[extracted_function_reduction.scala 659:35]
  assign br_24_clock = clock;
  assign br_24_reset = reset;
  assign br_24_io_enable_valid = bb_for_body15_lr_ph9_io_Out_3_valid; // @[extracted_function_reduction.scala 815:19]
  assign br_24_io_enable_bits_taskID = bb_for_body15_lr_ph9_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 815:19]
  assign br_24_io_enable_bits_control = bb_for_body15_lr_ph9_io_Out_3_bits_control; // @[extracted_function_reduction.scala 815:19]
  assign br_24_io_Out_0_ready = Loop_3_io_enable_ready; // @[extracted_function_reduction.scala 483:20]
  assign br_25_clock = clock;
  assign br_25_reset = reset;
  assign br_25_io_enable_valid = bb_for_cond_cleanup14_loopexit10_io_Out_0_valid; // @[extracted_function_reduction.scala 818:19]
  assign br_25_io_enable_bits_taskID = bb_for_cond_cleanup14_loopexit10_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 818:19]
  assign br_25_io_enable_bits_control = bb_for_cond_cleanup14_loopexit10_io_Out_0_bits_control; // @[extracted_function_reduction.scala 818:19]
  assign br_25_io_Out_0_ready = bb_for_cond_cleanup1411_io_predicateIn_0_ready; // @[extracted_function_reduction.scala 409:45]
  assign binaryOp_inc6126_clock = clock;
  assign binaryOp_inc6126_reset = reset;
  assign binaryOp_inc6126_io_enable_valid = bb_for_cond_cleanup1411_io_Out_1_valid; // @[extracted_function_reduction.scala 823:30]
  assign binaryOp_inc6126_io_enable_bits_taskID = bb_for_cond_cleanup1411_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 823:30]
  assign binaryOp_inc6126_io_enable_bits_control = bb_for_cond_cleanup1411_io_Out_1_bits_control; // @[extracted_function_reduction.scala 823:30]
  assign binaryOp_inc6126_io_Out_0_ready = Loop_4_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 709:29]
  assign binaryOp_inc6126_io_Out_1_ready = icmp_exitcond14727_io_LeftIO_ready; // @[extracted_function_reduction.scala 1098:32]
  assign binaryOp_inc6126_io_LeftIO_valid = phi_pw_conv_reduction_s1_y_014019_io_Out_2_valid; // @[extracted_function_reduction.scala 1092:30]
  assign binaryOp_inc6126_io_LeftIO_bits_data = phi_pw_conv_reduction_s1_y_014019_io_Out_2_bits_data; // @[extracted_function_reduction.scala 1092:30]
  assign binaryOp_inc6126_io_RightIO_valid = const1_io_Out_valid; // @[extracted_function_reduction.scala 1046:31]
  assign icmp_exitcond14727_clock = clock;
  assign icmp_exitcond14727_reset = reset;
  assign icmp_exitcond14727_io_enable_valid = bb_for_cond_cleanup1411_io_Out_2_valid; // @[extracted_function_reduction.scala 826:32]
  assign icmp_exitcond14727_io_enable_bits_taskID = bb_for_cond_cleanup1411_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 826:32]
  assign icmp_exitcond14727_io_enable_bits_control = bb_for_cond_cleanup1411_io_Out_2_bits_control; // @[extracted_function_reduction.scala 826:32]
  assign icmp_exitcond14727_io_Out_0_ready = br_28_io_CmpIO_ready; // @[extracted_function_reduction.scala 1100:18]
  assign icmp_exitcond14727_io_LeftIO_valid = binaryOp_inc6126_io_Out_1_valid; // @[extracted_function_reduction.scala 1098:32]
  assign icmp_exitcond14727_io_LeftIO_bits_data = binaryOp_inc6126_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1098:32]
  assign icmp_exitcond14727_io_RightIO_valid = Loop_4_io_OutLiveIn_field9_0_valid; // @[extracted_function_reduction.scala 653:33]
  assign icmp_exitcond14727_io_RightIO_bits_data = Loop_4_io_OutLiveIn_field9_0_bits_data; // @[extracted_function_reduction.scala 653:33]
  assign br_28_clock = clock;
  assign br_28_reset = reset;
  assign br_28_io_enable_valid = bb_for_cond_cleanup1411_io_Out_3_valid; // @[extracted_function_reduction.scala 829:19]
  assign br_28_io_enable_bits_taskID = bb_for_cond_cleanup1411_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 829:19]
  assign br_28_io_enable_bits_control = bb_for_cond_cleanup1411_io_Out_3_bits_control; // @[extracted_function_reduction.scala 829:19]
  assign br_28_io_CmpIO_valid = icmp_exitcond14727_io_Out_0_valid; // @[extracted_function_reduction.scala 1100:18]
  assign br_28_io_CmpIO_bits_taskID = icmp_exitcond14727_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 1100:18]
  assign br_28_io_CmpIO_bits_data = icmp_exitcond14727_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1100:18]
  assign br_28_io_TrueOutput_0_ready = Loop_4_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 493:27]
  assign br_28_io_FalseOutput_0_ready = Loop_4_io_loopBack_0_ready; // @[extracted_function_reduction.scala 491:25]
  assign phi_pw_conv_reduction_s1_x_013829_clock = clock;
  assign phi_pw_conv_reduction_s1_x_013829_reset = reset;
  assign phi_pw_conv_reduction_s1_x_013829_io_enable_valid = bb_for_body1512_io_Out_0_valid; // @[extracted_function_reduction.scala 832:47]
  assign phi_pw_conv_reduction_s1_x_013829_io_enable_bits_control = bb_for_body1512_io_Out_0_bits_control; // @[extracted_function_reduction.scala 832:47]
  assign phi_pw_conv_reduction_s1_x_013829_io_InData_0_valid = Loop_3_io_OutLiveIn_field8_0_valid; // @[extracted_function_reduction.scala 645:50]
  assign phi_pw_conv_reduction_s1_x_013829_io_InData_0_bits_taskID = Loop_3_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_reduction.scala 645:50]
  assign phi_pw_conv_reduction_s1_x_013829_io_InData_0_bits_data = Loop_3_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_reduction.scala 645:50]
  assign phi_pw_conv_reduction_s1_x_013829_io_InData_1_valid = Loop_3_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 729:50]
  assign phi_pw_conv_reduction_s1_x_013829_io_InData_1_bits_taskID = Loop_3_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 729:50]
  assign phi_pw_conv_reduction_s1_x_013829_io_InData_1_bits_data = Loop_3_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 729:50]
  assign phi_pw_conv_reduction_s1_x_013829_io_Mask_valid = bb_for_body1512_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 992:45]
  assign phi_pw_conv_reduction_s1_x_013829_io_Mask_bits = bb_for_body1512_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 992:45]
  assign phi_pw_conv_reduction_s1_x_013829_io_Out_0_ready = binaryOp_sub1630_io_LeftIO_ready; // @[extracted_function_reduction.scala 1102:30]
  assign phi_pw_conv_reduction_s1_x_013829_io_Out_1_ready = binaryOp_add1031_io_LeftIO_ready; // @[extracted_function_reduction.scala 1104:30]
  assign phi_pw_conv_reduction_s1_x_013829_io_Out_2_ready = binaryOp_inc5835_io_LeftIO_ready; // @[extracted_function_reduction.scala 1106:30]
  assign binaryOp_sub1630_clock = clock;
  assign binaryOp_sub1630_reset = reset;
  assign binaryOp_sub1630_io_enable_valid = bb_for_body1512_io_Out_1_valid; // @[extracted_function_reduction.scala 835:30]
  assign binaryOp_sub1630_io_enable_bits_taskID = bb_for_body1512_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 835:30]
  assign binaryOp_sub1630_io_enable_bits_control = bb_for_body1512_io_Out_1_bits_control; // @[extracted_function_reduction.scala 835:30]
  assign binaryOp_sub1630_io_Out_0_ready = Loop_2_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 527:25]
  assign binaryOp_sub1630_io_LeftIO_valid = phi_pw_conv_reduction_s1_x_013829_io_Out_0_valid; // @[extracted_function_reduction.scala 1102:30]
  assign binaryOp_sub1630_io_LeftIO_bits_data = phi_pw_conv_reduction_s1_x_013829_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1102:30]
  assign binaryOp_sub1630_io_RightIO_valid = Loop_3_io_OutLiveIn_field7_0_valid; // @[extracted_function_reduction.scala 643:31]
  assign binaryOp_sub1630_io_RightIO_bits_data = Loop_3_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_reduction.scala 643:31]
  assign binaryOp_add1031_clock = clock;
  assign binaryOp_add1031_reset = reset;
  assign binaryOp_add1031_io_enable_valid = bb_for_body1512_io_Out_2_valid; // @[extracted_function_reduction.scala 838:30]
  assign binaryOp_add1031_io_enable_bits_taskID = bb_for_body1512_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 838:30]
  assign binaryOp_add1031_io_enable_bits_control = bb_for_body1512_io_Out_2_bits_control; // @[extracted_function_reduction.scala 838:30]
  assign binaryOp_add1031_io_Out_0_ready = binaryOp_add1732_io_LeftIO_ready; // @[extracted_function_reduction.scala 1108:30]
  assign binaryOp_add1031_io_LeftIO_valid = phi_pw_conv_reduction_s1_x_013829_io_Out_1_valid; // @[extracted_function_reduction.scala 1104:30]
  assign binaryOp_add1031_io_LeftIO_bits_data = phi_pw_conv_reduction_s1_x_013829_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1104:30]
  assign binaryOp_add1031_io_RightIO_valid = Loop_3_io_OutLiveIn_field8_1_valid; // @[extracted_function_reduction.scala 647:31]
  assign binaryOp_add1031_io_RightIO_bits_data = Loop_3_io_OutLiveIn_field8_1_bits_data; // @[extracted_function_reduction.scala 647:31]
  assign binaryOp_add1732_clock = clock;
  assign binaryOp_add1732_reset = reset;
  assign binaryOp_add1732_io_enable_valid = bb_for_body1512_io_Out_3_valid; // @[extracted_function_reduction.scala 841:30]
  assign binaryOp_add1732_io_enable_bits_taskID = bb_for_body1512_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 841:30]
  assign binaryOp_add1732_io_enable_bits_control = bb_for_body1512_io_Out_3_bits_control; // @[extracted_function_reduction.scala 841:30]
  assign binaryOp_add1732_io_Out_0_ready = Gep_arrayidx5033_io_idx_0_ready; // @[extracted_function_reduction.scala 1110:30]
  assign binaryOp_add1732_io_LeftIO_valid = binaryOp_add1031_io_Out_0_valid; // @[extracted_function_reduction.scala 1108:30]
  assign binaryOp_add1732_io_LeftIO_bits_data = binaryOp_add1031_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1108:30]
  assign binaryOp_add1732_io_RightIO_valid = Loop_3_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 637:31]
  assign binaryOp_add1732_io_RightIO_bits_data = Loop_3_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 637:31]
  assign Gep_arrayidx5033_clock = clock;
  assign Gep_arrayidx5033_reset = reset;
  assign Gep_arrayidx5033_io_enable_valid = bb_for_body1512_io_Out_4_valid; // @[extracted_function_reduction.scala 844:30]
  assign Gep_arrayidx5033_io_enable_bits_taskID = bb_for_body1512_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 844:30]
  assign Gep_arrayidx5033_io_enable_bits_control = bb_for_body1512_io_Out_4_bits_control; // @[extracted_function_reduction.scala 844:30]
  assign Gep_arrayidx5033_io_Out_0_ready = Loop_2_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 529:25]
  assign Gep_arrayidx5033_io_baseAddress_valid = Loop_3_io_OutLiveIn_field5_0_valid; // @[extracted_function_reduction.scala 639:35]
  assign Gep_arrayidx5033_io_baseAddress_bits_taskID = Loop_3_io_OutLiveIn_field5_0_bits_taskID; // @[extracted_function_reduction.scala 639:35]
  assign Gep_arrayidx5033_io_baseAddress_bits_data = Loop_3_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_reduction.scala 639:35]
  assign Gep_arrayidx5033_io_idx_0_valid = binaryOp_add1732_io_Out_0_valid; // @[extracted_function_reduction.scala 1110:30]
  assign Gep_arrayidx5033_io_idx_0_bits_data = binaryOp_add1732_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1110:30]
  assign br_34_clock = clock;
  assign br_34_reset = reset;
  assign br_34_io_enable_valid = bb_for_body1512_io_Out_5_valid; // @[extracted_function_reduction.scala 847:19]
  assign br_34_io_enable_bits_taskID = bb_for_body1512_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 847:19]
  assign br_34_io_enable_bits_control = bb_for_body1512_io_Out_5_bits_control; // @[extracted_function_reduction.scala 847:19]
  assign br_34_io_Out_0_ready = Loop_2_io_enable_ready; // @[extracted_function_reduction.scala 477:20]
  assign binaryOp_inc5835_clock = clock;
  assign binaryOp_inc5835_reset = reset;
  assign binaryOp_inc5835_io_enable_valid = bb_for_cond_cleanup2013_io_Out_1_valid; // @[extracted_function_reduction.scala 852:30]
  assign binaryOp_inc5835_io_enable_bits_taskID = bb_for_cond_cleanup2013_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 852:30]
  assign binaryOp_inc5835_io_enable_bits_control = bb_for_cond_cleanup2013_io_Out_1_bits_control; // @[extracted_function_reduction.scala 852:30]
  assign binaryOp_inc5835_io_Out_0_ready = Loop_3_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 707:29]
  assign binaryOp_inc5835_io_Out_1_ready = icmp_exitcond14636_io_LeftIO_ready; // @[extracted_function_reduction.scala 1112:32]
  assign binaryOp_inc5835_io_LeftIO_valid = phi_pw_conv_reduction_s1_x_013829_io_Out_2_valid; // @[extracted_function_reduction.scala 1106:30]
  assign binaryOp_inc5835_io_LeftIO_bits_data = phi_pw_conv_reduction_s1_x_013829_io_Out_2_bits_data; // @[extracted_function_reduction.scala 1106:30]
  assign binaryOp_inc5835_io_RightIO_valid = const2_io_Out_valid; // @[extracted_function_reduction.scala 1048:31]
  assign icmp_exitcond14636_clock = clock;
  assign icmp_exitcond14636_reset = reset;
  assign icmp_exitcond14636_io_enable_valid = bb_for_cond_cleanup2013_io_Out_2_valid; // @[extracted_function_reduction.scala 855:32]
  assign icmp_exitcond14636_io_enable_bits_taskID = bb_for_cond_cleanup2013_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 855:32]
  assign icmp_exitcond14636_io_enable_bits_control = bb_for_cond_cleanup2013_io_Out_2_bits_control; // @[extracted_function_reduction.scala 855:32]
  assign icmp_exitcond14636_io_Out_0_ready = br_37_io_CmpIO_ready; // @[extracted_function_reduction.scala 1114:18]
  assign icmp_exitcond14636_io_LeftIO_valid = binaryOp_inc5835_io_Out_1_valid; // @[extracted_function_reduction.scala 1112:32]
  assign icmp_exitcond14636_io_LeftIO_bits_data = binaryOp_inc5835_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1112:32]
  assign icmp_exitcond14636_io_RightIO_valid = Loop_3_io_OutLiveIn_field6_0_valid; // @[extracted_function_reduction.scala 641:33]
  assign icmp_exitcond14636_io_RightIO_bits_data = Loop_3_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_reduction.scala 641:33]
  assign br_37_clock = clock;
  assign br_37_reset = reset;
  assign br_37_io_enable_valid = bb_for_cond_cleanup2013_io_Out_3_valid; // @[extracted_function_reduction.scala 858:19]
  assign br_37_io_enable_bits_taskID = bb_for_cond_cleanup2013_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 858:19]
  assign br_37_io_enable_bits_control = bb_for_cond_cleanup2013_io_Out_3_bits_control; // @[extracted_function_reduction.scala 858:19]
  assign br_37_io_CmpIO_valid = icmp_exitcond14636_io_Out_0_valid; // @[extracted_function_reduction.scala 1114:18]
  assign br_37_io_CmpIO_bits_taskID = icmp_exitcond14636_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 1114:18]
  assign br_37_io_CmpIO_bits_data = icmp_exitcond14636_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1114:18]
  assign br_37_io_TrueOutput_0_ready = Loop_3_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 487:27]
  assign br_37_io_FalseOutput_0_ready = Loop_3_io_loopBack_0_ready; // @[extracted_function_reduction.scala 485:25]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_clock = clock;
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_reset = reset;
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_enable_valid = bb_for_body2114_io_Out_1_valid; // @[extracted_function_reduction.scala 863:53]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_enable_bits_control = bb_for_body2114_io_Out_1_bits_control; // @[extracted_function_reduction.scala 863:53]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_0_valid = const3_io_Out_valid; // @[extracted_function_reduction.scala 1050:56]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_0_bits_taskID = const3_io_Out_bits_taskID; // @[extracted_function_reduction.scala 1050:56]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_valid = Loop_2_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 727:56]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_bits_taskID = Loop_2_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 727:56]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_1_bits_data = Loop_2_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 727:56]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_Mask_valid = bb_for_body2114_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 994:51]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_Mask_bits = bb_for_body2114_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 994:51]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_0_ready = binaryOp_mul2239_io_LeftIO_ready; // @[extracted_function_reduction.scala 1116:30]
  assign phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_1_ready = binaryOp_inc5548_io_LeftIO_ready; // @[extracted_function_reduction.scala 1118:30]
  assign binaryOp_mul2239_clock = clock;
  assign binaryOp_mul2239_reset = reset;
  assign binaryOp_mul2239_io_enable_valid = bb_for_body2114_io_Out_2_valid; // @[extracted_function_reduction.scala 866:30]
  assign binaryOp_mul2239_io_enable_bits_taskID = bb_for_body2114_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 866:30]
  assign binaryOp_mul2239_io_enable_bits_control = bb_for_body2114_io_Out_2_bits_control; // @[extracted_function_reduction.scala 866:30]
  assign binaryOp_mul2239_io_Out_0_ready = binaryOp_add2340_io_RightIO_ready; // @[extracted_function_reduction.scala 1120:31]
  assign binaryOp_mul2239_io_LeftIO_valid = phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_0_valid; // @[extracted_function_reduction.scala 1116:30]
  assign binaryOp_mul2239_io_LeftIO_bits_data = phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1116:30]
  assign binaryOp_mul2239_io_RightIO_valid = Loop_2_io_OutLiveIn_field5_0_valid; // @[extracted_function_reduction.scala 635:31]
  assign binaryOp_mul2239_io_RightIO_bits_data = Loop_2_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_reduction.scala 635:31]
  assign binaryOp_add2340_clock = clock;
  assign binaryOp_add2340_reset = reset;
  assign binaryOp_add2340_io_enable_valid = bb_for_body2114_io_Out_3_valid; // @[extracted_function_reduction.scala 869:30]
  assign binaryOp_add2340_io_enable_bits_taskID = bb_for_body2114_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 869:30]
  assign binaryOp_add2340_io_enable_bits_control = bb_for_body2114_io_Out_3_bits_control; // @[extracted_function_reduction.scala 869:30]
  assign binaryOp_add2340_io_Out_0_ready = Loop_1_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 519:25]
  assign binaryOp_add2340_io_LeftIO_valid = Loop_2_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 629:30]
  assign binaryOp_add2340_io_LeftIO_bits_data = Loop_2_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 629:30]
  assign binaryOp_add2340_io_RightIO_valid = binaryOp_mul2239_io_Out_0_valid; // @[extracted_function_reduction.scala 1120:31]
  assign binaryOp_add2340_io_RightIO_bits_data = binaryOp_mul2239_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1120:31]
  assign br_41_clock = clock;
  assign br_41_reset = reset;
  assign br_41_io_enable_valid = bb_for_body2114_io_Out_4_valid; // @[extracted_function_reduction.scala 872:19]
  assign br_41_io_enable_bits_taskID = bb_for_body2114_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 872:19]
  assign br_41_io_enable_bits_control = bb_for_body2114_io_Out_4_bits_control; // @[extracted_function_reduction.scala 872:19]
  assign br_41_io_Out_0_ready = Loop_1_io_enable_ready; // @[extracted_function_reduction.scala 471:20]
  assign phiadd38_lcssa_lcssa42_clock = clock;
  assign phiadd38_lcssa_lcssa42_reset = reset;
  assign phiadd38_lcssa_lcssa42_io_enable_valid = bb_for_cond_cleanup2615_io_Out_3_valid; // @[extracted_function_reduction.scala 881:36]
  assign phiadd38_lcssa_lcssa42_io_enable_bits_control = bb_for_cond_cleanup2615_io_Out_3_bits_control; // @[extracted_function_reduction.scala 881:36]
  assign phiadd38_lcssa_lcssa42_io_InData_0_valid = Loop_1_io_OutLiveOut_field0_0_valid; // @[extracted_function_reduction.scala 689:39]
  assign phiadd38_lcssa_lcssa42_io_InData_0_bits_taskID = Loop_1_io_OutLiveOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 689:39]
  assign phiadd38_lcssa_lcssa42_io_InData_0_bits_data = Loop_1_io_OutLiveOut_field0_0_bits_data; // @[extracted_function_reduction.scala 689:39]
  assign phiadd38_lcssa_lcssa42_io_Out_0_ready = binaryOp_mul4443_io_LeftIO_ready; // @[extracted_function_reduction.scala 1122:30]
  assign binaryOp_mul4443_clock = clock;
  assign binaryOp_mul4443_reset = reset;
  assign binaryOp_mul4443_io_enable_valid = bb_for_cond_cleanup2615_io_Out_4_valid; // @[extracted_function_reduction.scala 884:30]
  assign binaryOp_mul4443_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 884:30]
  assign binaryOp_mul4443_io_enable_bits_control = bb_for_cond_cleanup2615_io_Out_4_bits_control; // @[extracted_function_reduction.scala 884:30]
  assign binaryOp_mul4443_io_Out_0_ready = sextconv4744_io_Input_ready; // @[extracted_function_reduction.scala 1124:25]
  assign binaryOp_mul4443_io_LeftIO_valid = phiadd38_lcssa_lcssa42_io_Out_0_valid; // @[extracted_function_reduction.scala 1122:30]
  assign binaryOp_mul4443_io_LeftIO_bits_data = phiadd38_lcssa_lcssa42_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1122:30]
  assign binaryOp_mul4443_io_RightIO_valid = const4_io_Out_valid; // @[extracted_function_reduction.scala 1052:31]
  assign sextconv4744_clock = clock;
  assign sextconv4744_reset = reset;
  assign sextconv4744_io_Input_valid = binaryOp_mul4443_io_Out_0_valid; // @[extracted_function_reduction.scala 1124:25]
  assign sextconv4744_io_Input_bits_data = binaryOp_mul4443_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1124:25]
  assign sextconv4744_io_enable_valid = bb_for_cond_cleanup2615_io_Out_5_valid; // @[extracted_function_reduction.scala 887:26]
  assign sextconv4744_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 887:26]
  assign sextconv4744_io_Out_0_ready = binaryOp_add5246_io_RightIO_ready; // @[extracted_function_reduction.scala 1126:31]
  assign ld_45_clock = clock;
  assign ld_45_reset = reset;
  assign ld_45_io_enable_valid = bb_for_cond_cleanup2615_io_Out_6_valid; // @[extracted_function_reduction.scala 890:19]
  assign ld_45_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_6_bits_taskID; // @[extracted_function_reduction.scala 890:19]
  assign ld_45_io_enable_bits_control = bb_for_cond_cleanup2615_io_Out_6_bits_control; // @[extracted_function_reduction.scala 890:19]
  assign ld_45_io_Out_0_ready = binaryOp_add5246_io_LeftIO_ready; // @[extracted_function_reduction.scala 1128:30]
  assign ld_45_io_GepAddr_valid = Loop_2_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 631:20]
  assign ld_45_io_GepAddr_bits_predicate = Loop_2_io_OutLiveIn_field1_0_bits_predicate; // @[extracted_function_reduction.scala 631:20]
  assign ld_45_io_GepAddr_bits_taskID = Loop_2_io_OutLiveIn_field1_0_bits_taskID; // @[extracted_function_reduction.scala 631:20]
  assign ld_45_io_GepAddr_bits_data = Loop_2_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 631:20]
  assign ld_45_io_memReq_ready = MemCtrl_io_ReadIn_0_ready; // @[extracted_function_reduction.scala 1020:24]
  assign ld_45_io_memResp_valid = MemCtrl_io_ReadOut_0_valid; // @[extracted_function_reduction.scala 1022:20]
  assign ld_45_io_memResp_data = MemCtrl_io_ReadOut_0_data; // @[extracted_function_reduction.scala 1022:20]
  assign binaryOp_add5246_clock = clock;
  assign binaryOp_add5246_reset = reset;
  assign binaryOp_add5246_io_enable_valid = bb_for_cond_cleanup2615_io_Out_7_valid; // @[extracted_function_reduction.scala 893:30]
  assign binaryOp_add5246_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_7_bits_taskID; // @[extracted_function_reduction.scala 893:30]
  assign binaryOp_add5246_io_enable_bits_control = bb_for_cond_cleanup2615_io_Out_7_bits_control; // @[extracted_function_reduction.scala 893:30]
  assign binaryOp_add5246_io_Out_0_ready = st_47_io_inData_ready; // @[extracted_function_reduction.scala 1130:19]
  assign binaryOp_add5246_io_LeftIO_valid = ld_45_io_Out_0_valid; // @[extracted_function_reduction.scala 1128:30]
  assign binaryOp_add5246_io_LeftIO_bits_data = ld_45_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1128:30]
  assign binaryOp_add5246_io_RightIO_valid = sextconv4744_io_Out_0_valid; // @[extracted_function_reduction.scala 1126:31]
  assign binaryOp_add5246_io_RightIO_bits_data = sextconv4744_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1126:31]
  assign st_47_clock = clock;
  assign st_47_reset = reset;
  assign st_47_io_enable_valid = bb_for_cond_cleanup2615_io_Out_8_valid; // @[extracted_function_reduction.scala 896:19]
  assign st_47_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_8_bits_taskID; // @[extracted_function_reduction.scala 896:19]
  assign st_47_io_enable_bits_control = bb_for_cond_cleanup2615_io_Out_8_bits_control; // @[extracted_function_reduction.scala 896:19]
  assign st_47_io_GepAddr_valid = Loop_2_io_OutLiveIn_field1_1_valid; // @[extracted_function_reduction.scala 633:20]
  assign st_47_io_GepAddr_bits_taskID = Loop_2_io_OutLiveIn_field1_1_bits_taskID; // @[extracted_function_reduction.scala 633:20]
  assign st_47_io_GepAddr_bits_data = Loop_2_io_OutLiveIn_field1_1_bits_data; // @[extracted_function_reduction.scala 633:20]
  assign st_47_io_inData_valid = binaryOp_add5246_io_Out_0_valid; // @[extracted_function_reduction.scala 1130:19]
  assign st_47_io_inData_bits_taskID = binaryOp_add5246_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 1130:19]
  assign st_47_io_inData_bits_data = binaryOp_add5246_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1130:19]
  assign st_47_io_memReq_ready = MemCtrl_io_WriteIn_0_ready; // @[extracted_function_reduction.scala 1024:25]
  assign st_47_io_memResp_valid = MemCtrl_io_WriteOut_0_valid; // @[extracted_function_reduction.scala 1026:20]
  assign binaryOp_inc5548_clock = clock;
  assign binaryOp_inc5548_reset = reset;
  assign binaryOp_inc5548_io_enable_valid = bb_for_cond_cleanup2615_io_Out_9_valid; // @[extracted_function_reduction.scala 899:30]
  assign binaryOp_inc5548_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_9_bits_taskID; // @[extracted_function_reduction.scala 899:30]
  assign binaryOp_inc5548_io_enable_bits_control = bb_for_cond_cleanup2615_io_Out_9_bits_control; // @[extracted_function_reduction.scala 899:30]
  assign binaryOp_inc5548_io_Out_0_ready = Loop_2_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 705:29]
  assign binaryOp_inc5548_io_Out_1_ready = icmp_exitcond14549_io_LeftIO_ready; // @[extracted_function_reduction.scala 1132:32]
  assign binaryOp_inc5548_io_LeftIO_valid = phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_1_valid; // @[extracted_function_reduction.scala 1118:30]
  assign binaryOp_inc5548_io_LeftIO_bits_data = phi_pw_conv_reduction_s1_r_pw__x_013638_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1118:30]
  assign binaryOp_inc5548_io_RightIO_valid = const5_io_Out_valid; // @[extracted_function_reduction.scala 1054:31]
  assign icmp_exitcond14549_clock = clock;
  assign icmp_exitcond14549_reset = reset;
  assign icmp_exitcond14549_io_enable_valid = bb_for_cond_cleanup2615_io_Out_10_valid; // @[extracted_function_reduction.scala 902:32]
  assign icmp_exitcond14549_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_10_bits_taskID; // @[extracted_function_reduction.scala 902:32]
  assign icmp_exitcond14549_io_enable_bits_control = bb_for_cond_cleanup2615_io_Out_10_bits_control; // @[extracted_function_reduction.scala 902:32]
  assign icmp_exitcond14549_io_Out_0_ready = br_50_io_CmpIO_ready; // @[extracted_function_reduction.scala 1134:18]
  assign icmp_exitcond14549_io_LeftIO_valid = binaryOp_inc5548_io_Out_1_valid; // @[extracted_function_reduction.scala 1132:32]
  assign icmp_exitcond14549_io_LeftIO_bits_data = binaryOp_inc5548_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1132:32]
  assign icmp_exitcond14549_io_RightIO_valid = const6_io_Out_valid; // @[extracted_function_reduction.scala 1056:33]
  assign br_50_clock = clock;
  assign br_50_reset = reset;
  assign br_50_io_enable_valid = bb_for_cond_cleanup2615_io_Out_11_valid; // @[extracted_function_reduction.scala 905:19]
  assign br_50_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_11_bits_taskID; // @[extracted_function_reduction.scala 905:19]
  assign br_50_io_enable_bits_control = bb_for_cond_cleanup2615_io_Out_11_bits_control; // @[extracted_function_reduction.scala 905:19]
  assign br_50_io_CmpIO_valid = icmp_exitcond14549_io_Out_0_valid; // @[extracted_function_reduction.scala 1134:18]
  assign br_50_io_CmpIO_bits_taskID = icmp_exitcond14549_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 1134:18]
  assign br_50_io_CmpIO_bits_data = icmp_exitcond14549_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1134:18]
  assign br_50_io_TrueOutput_0_ready = Loop_2_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 481:27]
  assign br_50_io_FalseOutput_0_ready = Loop_2_io_loopBack_0_ready; // @[extracted_function_reduction.scala 479:25]
  assign phi_dw_conv_013551_clock = clock;
  assign phi_dw_conv_013551_reset = reset;
  assign phi_dw_conv_013551_io_enable_valid = bb_for_body2716_io_Out_2_valid; // @[extracted_function_reduction.scala 912:32]
  assign phi_dw_conv_013551_io_enable_bits_taskID = bb_for_body2716_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 912:32]
  assign phi_dw_conv_013551_io_enable_bits_control = bb_for_body2716_io_Out_2_bits_control; // @[extracted_function_reduction.scala 912:32]
  assign phi_dw_conv_013551_io_InData_0_valid = const7_io_Out_valid; // @[extracted_function_reduction.scala 1058:35]
  assign phi_dw_conv_013551_io_InData_0_bits_taskID = const7_io_Out_bits_taskID; // @[extracted_function_reduction.scala 1058:35]
  assign phi_dw_conv_013551_io_InData_1_valid = Loop_1_io_CarryDepenOut_field1_0_valid; // @[extracted_function_reduction.scala 725:35]
  assign phi_dw_conv_013551_io_InData_1_bits_taskID = Loop_1_io_CarryDepenOut_field1_0_bits_taskID; // @[extracted_function_reduction.scala 725:35]
  assign phi_dw_conv_013551_io_InData_1_bits_data = Loop_1_io_CarryDepenOut_field1_0_bits_data; // @[extracted_function_reduction.scala 725:35]
  assign phi_dw_conv_013551_io_Mask_valid = bb_for_body2716_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 998:30]
  assign phi_dw_conv_013551_io_Mask_bits = bb_for_body2716_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 998:30]
  assign phi_dw_conv_013551_io_Out_0_ready = Loop_0_io_InLiveIn_0_ready; // @[extracted_function_reduction.scala 513:25]
  assign phi_dw_conv_s1_r_dw__y_013452_clock = clock;
  assign phi_dw_conv_s1_r_dw__y_013452_reset = reset;
  assign phi_dw_conv_s1_r_dw__y_013452_io_enable_valid = bb_for_body2716_io_Out_3_valid; // @[extracted_function_reduction.scala 915:43]
  assign phi_dw_conv_s1_r_dw__y_013452_io_enable_bits_control = bb_for_body2716_io_Out_3_bits_control; // @[extracted_function_reduction.scala 915:43]
  assign phi_dw_conv_s1_r_dw__y_013452_io_InData_0_valid = const8_io_Out_valid; // @[extracted_function_reduction.scala 1060:46]
  assign phi_dw_conv_s1_r_dw__y_013452_io_InData_0_bits_taskID = const8_io_Out_bits_taskID; // @[extracted_function_reduction.scala 1060:46]
  assign phi_dw_conv_s1_r_dw__y_013452_io_InData_1_valid = Loop_1_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 723:46]
  assign phi_dw_conv_s1_r_dw__y_013452_io_InData_1_bits_taskID = Loop_1_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 723:46]
  assign phi_dw_conv_s1_r_dw__y_013452_io_InData_1_bits_data = Loop_1_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 723:46]
  assign phi_dw_conv_s1_r_dw__y_013452_io_Mask_valid = bb_for_body2716_io_MaskBB_1_valid; // @[extracted_function_reduction.scala 1000:41]
  assign phi_dw_conv_s1_r_dw__y_013452_io_Mask_bits = bb_for_body2716_io_MaskBB_1_bits; // @[extracted_function_reduction.scala 1000:41]
  assign phi_dw_conv_s1_r_dw__y_013452_io_Out_0_ready = binaryOp_add2853_io_LeftIO_ready; // @[extracted_function_reduction.scala 1136:30]
  assign phi_dw_conv_s1_r_dw__y_013452_io_Out_1_ready = binaryOp_inc4158_io_LeftIO_ready; // @[extracted_function_reduction.scala 1138:30]
  assign binaryOp_add2853_clock = clock;
  assign binaryOp_add2853_reset = reset;
  assign binaryOp_add2853_io_enable_valid = bb_for_body2716_io_Out_4_valid; // @[extracted_function_reduction.scala 918:30]
  assign binaryOp_add2853_io_enable_bits_taskID = bb_for_body2716_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 918:30]
  assign binaryOp_add2853_io_enable_bits_control = bb_for_body2716_io_Out_4_bits_control; // @[extracted_function_reduction.scala 918:30]
  assign binaryOp_add2853_io_Out_0_ready = binaryOp_mul2954_io_LeftIO_ready; // @[extracted_function_reduction.scala 1140:30]
  assign binaryOp_add2853_io_LeftIO_valid = phi_dw_conv_s1_r_dw__y_013452_io_Out_0_valid; // @[extracted_function_reduction.scala 1136:30]
  assign binaryOp_add2853_io_LeftIO_bits_data = phi_dw_conv_s1_r_dw__y_013452_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1136:30]
  assign binaryOp_add2853_io_RightIO_valid = Loop_1_io_OutLiveIn_field3_0_valid; // @[extracted_function_reduction.scala 627:31]
  assign binaryOp_add2853_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_reduction.scala 627:31]
  assign binaryOp_mul2954_clock = clock;
  assign binaryOp_mul2954_reset = reset;
  assign binaryOp_mul2954_io_enable_valid = bb_for_body2716_io_Out_5_valid; // @[extracted_function_reduction.scala 921:30]
  assign binaryOp_mul2954_io_enable_bits_taskID = bb_for_body2716_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 921:30]
  assign binaryOp_mul2954_io_enable_bits_control = bb_for_body2716_io_Out_5_bits_control; // @[extracted_function_reduction.scala 921:30]
  assign binaryOp_mul2954_io_Out_0_ready = binaryOp_add3055_io_RightIO_ready; // @[extracted_function_reduction.scala 1142:31]
  assign binaryOp_mul2954_io_LeftIO_valid = binaryOp_add2853_io_Out_0_valid; // @[extracted_function_reduction.scala 1140:30]
  assign binaryOp_mul2954_io_LeftIO_bits_data = binaryOp_add2853_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1140:30]
  assign binaryOp_mul2954_io_RightIO_valid = Loop_1_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 625:31]
  assign binaryOp_mul2954_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 625:31]
  assign binaryOp_add3055_clock = clock;
  assign binaryOp_add3055_reset = reset;
  assign binaryOp_add3055_io_enable_valid = bb_for_body2716_io_Out_6_valid; // @[extracted_function_reduction.scala 924:30]
  assign binaryOp_add3055_io_enable_bits_taskID = bb_for_body2716_io_Out_6_bits_taskID; // @[extracted_function_reduction.scala 924:30]
  assign binaryOp_add3055_io_enable_bits_control = bb_for_body2716_io_Out_6_bits_control; // @[extracted_function_reduction.scala 924:30]
  assign binaryOp_add3055_io_Out_0_ready = Loop_0_io_InLiveIn_1_ready; // @[extracted_function_reduction.scala 515:25]
  assign binaryOp_add3055_io_LeftIO_valid = Loop_1_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 623:30]
  assign binaryOp_add3055_io_LeftIO_bits_data = Loop_1_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 623:30]
  assign binaryOp_add3055_io_RightIO_valid = binaryOp_mul2954_io_Out_0_valid; // @[extracted_function_reduction.scala 1142:31]
  assign binaryOp_add3055_io_RightIO_bits_data = binaryOp_mul2954_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1142:31]
  assign br_56_clock = clock;
  assign br_56_reset = reset;
  assign br_56_io_enable_valid = bb_for_body2716_io_Out_7_valid; // @[extracted_function_reduction.scala 927:19]
  assign br_56_io_enable_bits_taskID = bb_for_body2716_io_Out_7_bits_taskID; // @[extracted_function_reduction.scala 927:19]
  assign br_56_io_enable_bits_control = bb_for_body2716_io_Out_7_bits_control; // @[extracted_function_reduction.scala 927:19]
  assign br_56_io_Out_0_ready = Loop_0_io_enable_ready; // @[extracted_function_reduction.scala 465:20]
  assign phiadd38_lcssa57_clock = clock;
  assign phiadd38_lcssa57_reset = reset;
  assign phiadd38_lcssa57_io_enable_valid = bb_for_cond_cleanup3317_io_Out_2_valid; // @[extracted_function_reduction.scala 934:30]
  assign phiadd38_lcssa57_io_enable_bits_taskID = bb_for_cond_cleanup3317_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 934:30]
  assign phiadd38_lcssa57_io_enable_bits_control = bb_for_cond_cleanup3317_io_Out_2_bits_control; // @[extracted_function_reduction.scala 934:30]
  assign phiadd38_lcssa57_io_InData_0_valid = Loop_0_io_OutLiveOut_field0_0_valid; // @[extracted_function_reduction.scala 687:33]
  assign phiadd38_lcssa57_io_InData_0_bits_taskID = Loop_0_io_OutLiveOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 687:33]
  assign phiadd38_lcssa57_io_InData_0_bits_data = Loop_0_io_OutLiveOut_field0_0_bits_data; // @[extracted_function_reduction.scala 687:33]
  assign phiadd38_lcssa57_io_Out_0_ready = Loop_1_io_InLiveOut_0_ready; // @[extracted_function_reduction.scala 679:26]
  assign phiadd38_lcssa57_io_Out_1_ready = Loop_1_io_CarryDepenIn_1_ready; // @[extracted_function_reduction.scala 703:29]
  assign binaryOp_inc4158_clock = clock;
  assign binaryOp_inc4158_reset = reset;
  assign binaryOp_inc4158_io_enable_valid = bb_for_cond_cleanup3317_io_Out_3_valid; // @[extracted_function_reduction.scala 937:30]
  assign binaryOp_inc4158_io_enable_bits_taskID = bb_for_cond_cleanup3317_io_Out_3_bits_taskID; // @[extracted_function_reduction.scala 937:30]
  assign binaryOp_inc4158_io_enable_bits_control = bb_for_cond_cleanup3317_io_Out_3_bits_control; // @[extracted_function_reduction.scala 937:30]
  assign binaryOp_inc4158_io_Out_0_ready = Loop_1_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 701:29]
  assign binaryOp_inc4158_io_Out_1_ready = icmp_exitcond14459_io_LeftIO_ready; // @[extracted_function_reduction.scala 1144:32]
  assign binaryOp_inc4158_io_LeftIO_valid = phi_dw_conv_s1_r_dw__y_013452_io_Out_1_valid; // @[extracted_function_reduction.scala 1138:30]
  assign binaryOp_inc4158_io_LeftIO_bits_data = phi_dw_conv_s1_r_dw__y_013452_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1138:30]
  assign binaryOp_inc4158_io_RightIO_valid = const9_io_Out_valid; // @[extracted_function_reduction.scala 1062:31]
  assign icmp_exitcond14459_clock = clock;
  assign icmp_exitcond14459_reset = reset;
  assign icmp_exitcond14459_io_enable_valid = bb_for_cond_cleanup3317_io_Out_4_valid; // @[extracted_function_reduction.scala 940:32]
  assign icmp_exitcond14459_io_enable_bits_taskID = bb_for_cond_cleanup3317_io_Out_4_bits_taskID; // @[extracted_function_reduction.scala 940:32]
  assign icmp_exitcond14459_io_enable_bits_control = bb_for_cond_cleanup3317_io_Out_4_bits_control; // @[extracted_function_reduction.scala 940:32]
  assign icmp_exitcond14459_io_Out_0_ready = br_60_io_CmpIO_ready; // @[extracted_function_reduction.scala 1146:18]
  assign icmp_exitcond14459_io_LeftIO_valid = binaryOp_inc4158_io_Out_1_valid; // @[extracted_function_reduction.scala 1144:32]
  assign icmp_exitcond14459_io_LeftIO_bits_data = binaryOp_inc4158_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1144:32]
  assign icmp_exitcond14459_io_RightIO_valid = const10_io_Out_valid; // @[extracted_function_reduction.scala 1064:33]
  assign br_60_clock = clock;
  assign br_60_reset = reset;
  assign br_60_io_enable_valid = bb_for_cond_cleanup3317_io_Out_5_valid; // @[extracted_function_reduction.scala 943:19]
  assign br_60_io_enable_bits_taskID = bb_for_cond_cleanup3317_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 943:19]
  assign br_60_io_enable_bits_control = bb_for_cond_cleanup3317_io_Out_5_bits_control; // @[extracted_function_reduction.scala 943:19]
  assign br_60_io_CmpIO_valid = icmp_exitcond14459_io_Out_0_valid; // @[extracted_function_reduction.scala 1146:18]
  assign br_60_io_CmpIO_bits_taskID = icmp_exitcond14459_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 1146:18]
  assign br_60_io_CmpIO_bits_data = icmp_exitcond14459_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1146:18]
  assign br_60_io_TrueOutput_0_ready = Loop_1_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 475:27]
  assign br_60_io_FalseOutput_0_ready = Loop_1_io_loopBack_0_ready; // @[extracted_function_reduction.scala 473:25]
  assign phi_dw_conv_113361_clock = clock;
  assign phi_dw_conv_113361_reset = reset;
  assign phi_dw_conv_113361_io_enable_valid = bb_for_body3418_io_Out_3_valid; // @[extracted_function_reduction.scala 952:32]
  assign phi_dw_conv_113361_io_enable_bits_control = bb_for_body3418_io_Out_3_bits_control; // @[extracted_function_reduction.scala 952:32]
  assign phi_dw_conv_113361_io_InData_0_valid = Loop_0_io_OutLiveIn_field0_0_valid; // @[extracted_function_reduction.scala 617:35]
  assign phi_dw_conv_113361_io_InData_0_bits_taskID = Loop_0_io_OutLiveIn_field0_0_bits_taskID; // @[extracted_function_reduction.scala 617:35]
  assign phi_dw_conv_113361_io_InData_0_bits_data = Loop_0_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_reduction.scala 617:35]
  assign phi_dw_conv_113361_io_InData_1_valid = Loop_0_io_CarryDepenOut_field0_0_valid; // @[extracted_function_reduction.scala 719:35]
  assign phi_dw_conv_113361_io_InData_1_bits_taskID = Loop_0_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_reduction.scala 719:35]
  assign phi_dw_conv_113361_io_InData_1_bits_data = Loop_0_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_reduction.scala 719:35]
  assign phi_dw_conv_113361_io_Mask_valid = bb_for_body3418_io_MaskBB_0_valid; // @[extracted_function_reduction.scala 1004:30]
  assign phi_dw_conv_113361_io_Mask_bits = bb_for_body3418_io_MaskBB_0_bits; // @[extracted_function_reduction.scala 1004:30]
  assign phi_dw_conv_113361_io_Out_0_ready = binaryOp_add3867_io_LeftIO_ready; // @[extracted_function_reduction.scala 1148:30]
  assign phi_dw_conv_s1_r_dw__x_013262_clock = clock;
  assign phi_dw_conv_s1_r_dw__x_013262_reset = reset;
  assign phi_dw_conv_s1_r_dw__x_013262_io_enable_valid = bb_for_body3418_io_Out_4_valid; // @[extracted_function_reduction.scala 955:43]
  assign phi_dw_conv_s1_r_dw__x_013262_io_enable_bits_control = bb_for_body3418_io_Out_4_bits_control; // @[extracted_function_reduction.scala 955:43]
  assign phi_dw_conv_s1_r_dw__x_013262_io_InData_0_valid = const11_io_Out_valid; // @[extracted_function_reduction.scala 1066:46]
  assign phi_dw_conv_s1_r_dw__x_013262_io_InData_0_bits_taskID = const11_io_Out_bits_taskID; // @[extracted_function_reduction.scala 1066:46]
  assign phi_dw_conv_s1_r_dw__x_013262_io_InData_1_valid = Loop_0_io_CarryDepenOut_field1_0_valid; // @[extracted_function_reduction.scala 721:46]
  assign phi_dw_conv_s1_r_dw__x_013262_io_InData_1_bits_taskID = Loop_0_io_CarryDepenOut_field1_0_bits_taskID; // @[extracted_function_reduction.scala 721:46]
  assign phi_dw_conv_s1_r_dw__x_013262_io_InData_1_bits_data = Loop_0_io_CarryDepenOut_field1_0_bits_data; // @[extracted_function_reduction.scala 721:46]
  assign phi_dw_conv_s1_r_dw__x_013262_io_Mask_valid = bb_for_body3418_io_MaskBB_1_valid; // @[extracted_function_reduction.scala 1006:41]
  assign phi_dw_conv_s1_r_dw__x_013262_io_Mask_bits = bb_for_body3418_io_MaskBB_1_bits; // @[extracted_function_reduction.scala 1006:41]
  assign phi_dw_conv_s1_r_dw__x_013262_io_Out_0_ready = binaryOp_add3563_io_RightIO_ready; // @[extracted_function_reduction.scala 1150:31]
  assign phi_dw_conv_s1_r_dw__x_013262_io_Out_1_ready = binaryOp_inc68_io_LeftIO_ready; // @[extracted_function_reduction.scala 1152:28]
  assign binaryOp_add3563_clock = clock;
  assign binaryOp_add3563_reset = reset;
  assign binaryOp_add3563_io_enable_valid = bb_for_body3418_io_Out_5_valid; // @[extracted_function_reduction.scala 958:30]
  assign binaryOp_add3563_io_enable_bits_taskID = bb_for_body3418_io_Out_5_bits_taskID; // @[extracted_function_reduction.scala 958:30]
  assign binaryOp_add3563_io_enable_bits_control = bb_for_body3418_io_Out_5_bits_control; // @[extracted_function_reduction.scala 958:30]
  assign binaryOp_add3563_io_Out_0_ready = Gep_arrayidx64_io_idx_0_ready; // @[extracted_function_reduction.scala 1154:28]
  assign binaryOp_add3563_io_LeftIO_valid = Loop_0_io_OutLiveIn_field1_0_valid; // @[extracted_function_reduction.scala 619:30]
  assign binaryOp_add3563_io_LeftIO_bits_data = Loop_0_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_reduction.scala 619:30]
  assign binaryOp_add3563_io_RightIO_valid = phi_dw_conv_s1_r_dw__x_013262_io_Out_0_valid; // @[extracted_function_reduction.scala 1150:31]
  assign binaryOp_add3563_io_RightIO_bits_data = phi_dw_conv_s1_r_dw__x_013262_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1150:31]
  assign Gep_arrayidx64_clock = clock;
  assign Gep_arrayidx64_reset = reset;
  assign Gep_arrayidx64_io_enable_valid = bb_for_body3418_io_Out_6_valid; // @[extracted_function_reduction.scala 961:28]
  assign Gep_arrayidx64_io_enable_bits_taskID = bb_for_body3418_io_Out_6_bits_taskID; // @[extracted_function_reduction.scala 961:28]
  assign Gep_arrayidx64_io_enable_bits_control = bb_for_body3418_io_Out_6_bits_control; // @[extracted_function_reduction.scala 961:28]
  assign Gep_arrayidx64_io_Out_0_ready = ld_65_io_GepAddr_ready; // @[extracted_function_reduction.scala 1156:20]
  assign Gep_arrayidx64_io_baseAddress_valid = Loop_0_io_OutLiveIn_field2_0_valid; // @[extracted_function_reduction.scala 621:33]
  assign Gep_arrayidx64_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field2_0_bits_taskID; // @[extracted_function_reduction.scala 621:33]
  assign Gep_arrayidx64_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_reduction.scala 621:33]
  assign Gep_arrayidx64_io_idx_0_valid = binaryOp_add3563_io_Out_0_valid; // @[extracted_function_reduction.scala 1154:28]
  assign Gep_arrayidx64_io_idx_0_bits_data = binaryOp_add3563_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1154:28]
  assign ld_65_clock = clock;
  assign ld_65_reset = reset;
  assign ld_65_io_enable_valid = bb_for_body3418_io_Out_7_valid; // @[extracted_function_reduction.scala 964:19]
  assign ld_65_io_enable_bits_taskID = bb_for_body3418_io_Out_7_bits_taskID; // @[extracted_function_reduction.scala 964:19]
  assign ld_65_io_enable_bits_control = bb_for_body3418_io_Out_7_bits_control; // @[extracted_function_reduction.scala 964:19]
  assign ld_65_io_Out_0_ready = sextconv3766_io_Input_ready; // @[extracted_function_reduction.scala 1158:25]
  assign ld_65_io_GepAddr_valid = Gep_arrayidx64_io_Out_0_valid; // @[extracted_function_reduction.scala 1156:20]
  assign ld_65_io_GepAddr_bits_predicate = Gep_arrayidx64_io_Out_0_bits_predicate; // @[extracted_function_reduction.scala 1156:20]
  assign ld_65_io_GepAddr_bits_taskID = Gep_arrayidx64_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 1156:20]
  assign ld_65_io_GepAddr_bits_data = Gep_arrayidx64_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1156:20]
  assign ld_65_io_memReq_ready = MemCtrl_io_ReadIn_1_ready; // @[extracted_function_reduction.scala 1028:24]
  assign ld_65_io_memResp_valid = MemCtrl_io_ReadOut_1_valid; // @[extracted_function_reduction.scala 1030:20]
  assign ld_65_io_memResp_data = MemCtrl_io_ReadOut_1_data; // @[extracted_function_reduction.scala 1030:20]
  assign sextconv3766_clock = clock;
  assign sextconv3766_reset = reset;
  assign sextconv3766_io_Input_valid = ld_65_io_Out_0_valid; // @[extracted_function_reduction.scala 1158:25]
  assign sextconv3766_io_Input_bits_data = ld_65_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1158:25]
  assign sextconv3766_io_enable_valid = bb_for_body3418_io_Out_8_valid; // @[extracted_function_reduction.scala 967:26]
  assign sextconv3766_io_enable_bits_taskID = bb_for_body3418_io_Out_8_bits_taskID; // @[extracted_function_reduction.scala 967:26]
  assign sextconv3766_io_Out_0_ready = binaryOp_add3867_io_RightIO_ready; // @[extracted_function_reduction.scala 1160:31]
  assign binaryOp_add3867_clock = clock;
  assign binaryOp_add3867_reset = reset;
  assign binaryOp_add3867_io_enable_valid = bb_for_body3418_io_Out_9_valid; // @[extracted_function_reduction.scala 970:30]
  assign binaryOp_add3867_io_enable_bits_taskID = bb_for_body3418_io_Out_9_bits_taskID; // @[extracted_function_reduction.scala 970:30]
  assign binaryOp_add3867_io_enable_bits_control = bb_for_body3418_io_Out_9_bits_control; // @[extracted_function_reduction.scala 970:30]
  assign binaryOp_add3867_io_Out_0_ready = Loop_0_io_InLiveOut_0_ready; // @[extracted_function_reduction.scala 677:26]
  assign binaryOp_add3867_io_Out_1_ready = Loop_0_io_CarryDepenIn_0_ready; // @[extracted_function_reduction.scala 697:29]
  assign binaryOp_add3867_io_LeftIO_valid = phi_dw_conv_113361_io_Out_0_valid; // @[extracted_function_reduction.scala 1148:30]
  assign binaryOp_add3867_io_LeftIO_bits_data = phi_dw_conv_113361_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1148:30]
  assign binaryOp_add3867_io_RightIO_valid = sextconv3766_io_Out_0_valid; // @[extracted_function_reduction.scala 1160:31]
  assign binaryOp_add3867_io_RightIO_bits_data = sextconv3766_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1160:31]
  assign binaryOp_inc68_clock = clock;
  assign binaryOp_inc68_reset = reset;
  assign binaryOp_inc68_io_enable_valid = bb_for_body3418_io_Out_10_valid; // @[extracted_function_reduction.scala 973:28]
  assign binaryOp_inc68_io_enable_bits_taskID = bb_for_body3418_io_Out_10_bits_taskID; // @[extracted_function_reduction.scala 973:28]
  assign binaryOp_inc68_io_enable_bits_control = bb_for_body3418_io_Out_10_bits_control; // @[extracted_function_reduction.scala 973:28]
  assign binaryOp_inc68_io_Out_0_ready = Loop_0_io_CarryDepenIn_1_ready; // @[extracted_function_reduction.scala 699:29]
  assign binaryOp_inc68_io_Out_1_ready = icmp_exitcond69_io_LeftIO_ready; // @[extracted_function_reduction.scala 1162:29]
  assign binaryOp_inc68_io_LeftIO_valid = phi_dw_conv_s1_r_dw__x_013262_io_Out_1_valid; // @[extracted_function_reduction.scala 1152:28]
  assign binaryOp_inc68_io_LeftIO_bits_data = phi_dw_conv_s1_r_dw__x_013262_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1152:28]
  assign binaryOp_inc68_io_RightIO_valid = const12_io_Out_valid; // @[extracted_function_reduction.scala 1068:29]
  assign icmp_exitcond69_clock = clock;
  assign icmp_exitcond69_reset = reset;
  assign icmp_exitcond69_io_enable_valid = bb_for_body3418_io_Out_11_valid; // @[extracted_function_reduction.scala 976:29]
  assign icmp_exitcond69_io_enable_bits_taskID = bb_for_body3418_io_Out_11_bits_taskID; // @[extracted_function_reduction.scala 976:29]
  assign icmp_exitcond69_io_enable_bits_control = bb_for_body3418_io_Out_11_bits_control; // @[extracted_function_reduction.scala 976:29]
  assign icmp_exitcond69_io_Out_0_ready = br_70_io_CmpIO_ready; // @[extracted_function_reduction.scala 1164:18]
  assign icmp_exitcond69_io_LeftIO_valid = binaryOp_inc68_io_Out_1_valid; // @[extracted_function_reduction.scala 1162:29]
  assign icmp_exitcond69_io_LeftIO_bits_data = binaryOp_inc68_io_Out_1_bits_data; // @[extracted_function_reduction.scala 1162:29]
  assign icmp_exitcond69_io_RightIO_valid = const13_io_Out_valid; // @[extracted_function_reduction.scala 1070:30]
  assign br_70_clock = clock;
  assign br_70_reset = reset;
  assign br_70_io_enable_valid = bb_for_body3418_io_Out_12_valid; // @[extracted_function_reduction.scala 979:19]
  assign br_70_io_enable_bits_taskID = bb_for_body3418_io_Out_12_bits_taskID; // @[extracted_function_reduction.scala 979:19]
  assign br_70_io_enable_bits_control = bb_for_body3418_io_Out_12_bits_control; // @[extracted_function_reduction.scala 979:19]
  assign br_70_io_CmpIO_valid = icmp_exitcond69_io_Out_0_valid; // @[extracted_function_reduction.scala 1164:18]
  assign br_70_io_CmpIO_bits_taskID = icmp_exitcond69_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 1164:18]
  assign br_70_io_CmpIO_bits_data = icmp_exitcond69_io_Out_0_bits_data; // @[extracted_function_reduction.scala 1164:18]
  assign br_70_io_TrueOutput_0_ready = Loop_0_io_loopFinish_0_ready; // @[extracted_function_reduction.scala 469:27]
  assign br_70_io_FalseOutput_0_ready = Loop_0_io_loopBack_0_ready; // @[extracted_function_reduction.scala 467:25]
  assign const0_clock = clock;
  assign const0_reset = reset;
  assign const0_io_enable_valid = bb_for_cond_cleanup67_io_Out_0_valid; // @[extracted_function_reduction.scala 789:20]
  assign const0_io_enable_bits_taskID = bb_for_cond_cleanup67_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 789:20]
  assign const0_io_Out_ready = binaryOp_inc6416_io_RightIO_ready; // @[extracted_function_reduction.scala 1044:31]
  assign const1_clock = clock;
  assign const1_reset = reset;
  assign const1_io_enable_valid = bb_for_cond_cleanup1411_io_Out_0_valid; // @[extracted_function_reduction.scala 821:20]
  assign const1_io_enable_bits_taskID = bb_for_cond_cleanup1411_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 821:20]
  assign const1_io_Out_ready = binaryOp_inc6126_io_RightIO_ready; // @[extracted_function_reduction.scala 1046:31]
  assign const2_clock = clock;
  assign const2_reset = reset;
  assign const2_io_enable_valid = bb_for_cond_cleanup2013_io_Out_0_valid; // @[extracted_function_reduction.scala 850:20]
  assign const2_io_enable_bits_taskID = bb_for_cond_cleanup2013_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 850:20]
  assign const2_io_Out_ready = binaryOp_inc5835_io_RightIO_ready; // @[extracted_function_reduction.scala 1048:31]
  assign const3_clock = clock;
  assign const3_reset = reset;
  assign const3_io_enable_valid = bb_for_body2114_io_Out_0_valid; // @[extracted_function_reduction.scala 861:20]
  assign const3_io_enable_bits_taskID = bb_for_body2114_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 861:20]
  assign const3_io_Out_ready = phi_pw_conv_reduction_s1_r_pw__x_013638_io_InData_0_ready; // @[extracted_function_reduction.scala 1050:56]
  assign const4_clock = clock;
  assign const4_reset = reset;
  assign const4_io_enable_valid = bb_for_cond_cleanup2615_io_Out_0_valid; // @[extracted_function_reduction.scala 875:20]
  assign const4_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 875:20]
  assign const4_io_Out_ready = binaryOp_mul4443_io_RightIO_ready; // @[extracted_function_reduction.scala 1052:31]
  assign const5_clock = clock;
  assign const5_reset = reset;
  assign const5_io_enable_valid = bb_for_cond_cleanup2615_io_Out_1_valid; // @[extracted_function_reduction.scala 877:20]
  assign const5_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 877:20]
  assign const5_io_Out_ready = binaryOp_inc5548_io_RightIO_ready; // @[extracted_function_reduction.scala 1054:31]
  assign const6_clock = clock;
  assign const6_reset = reset;
  assign const6_io_enable_valid = bb_for_cond_cleanup2615_io_Out_2_valid; // @[extracted_function_reduction.scala 879:20]
  assign const6_io_enable_bits_taskID = bb_for_cond_cleanup2615_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 879:20]
  assign const6_io_Out_ready = icmp_exitcond14549_io_RightIO_ready; // @[extracted_function_reduction.scala 1056:33]
  assign const7_clock = clock;
  assign const7_reset = reset;
  assign const7_io_enable_valid = bb_for_body2716_io_Out_0_valid; // @[extracted_function_reduction.scala 908:20]
  assign const7_io_enable_bits_taskID = bb_for_body2716_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 908:20]
  assign const7_io_Out_ready = phi_dw_conv_013551_io_InData_0_ready; // @[extracted_function_reduction.scala 1058:35]
  assign const8_clock = clock;
  assign const8_reset = reset;
  assign const8_io_enable_valid = bb_for_body2716_io_Out_1_valid; // @[extracted_function_reduction.scala 910:20]
  assign const8_io_enable_bits_taskID = bb_for_body2716_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 910:20]
  assign const8_io_Out_ready = phi_dw_conv_s1_r_dw__y_013452_io_InData_0_ready; // @[extracted_function_reduction.scala 1060:46]
  assign const9_clock = clock;
  assign const9_reset = reset;
  assign const9_io_enable_valid = bb_for_cond_cleanup3317_io_Out_0_valid; // @[extracted_function_reduction.scala 930:20]
  assign const9_io_enable_bits_taskID = bb_for_cond_cleanup3317_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 930:20]
  assign const9_io_Out_ready = binaryOp_inc4158_io_RightIO_ready; // @[extracted_function_reduction.scala 1062:31]
  assign const10_clock = clock;
  assign const10_reset = reset;
  assign const10_io_enable_valid = bb_for_cond_cleanup3317_io_Out_1_valid; // @[extracted_function_reduction.scala 932:21]
  assign const10_io_enable_bits_taskID = bb_for_cond_cleanup3317_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 932:21]
  assign const10_io_Out_ready = icmp_exitcond14459_io_RightIO_ready; // @[extracted_function_reduction.scala 1064:33]
  assign const11_clock = clock;
  assign const11_reset = reset;
  assign const11_io_enable_valid = bb_for_body3418_io_Out_0_valid; // @[extracted_function_reduction.scala 946:21]
  assign const11_io_enable_bits_taskID = bb_for_body3418_io_Out_0_bits_taskID; // @[extracted_function_reduction.scala 946:21]
  assign const11_io_Out_ready = phi_dw_conv_s1_r_dw__x_013262_io_InData_0_ready; // @[extracted_function_reduction.scala 1066:46]
  assign const12_clock = clock;
  assign const12_reset = reset;
  assign const12_io_enable_valid = bb_for_body3418_io_Out_1_valid; // @[extracted_function_reduction.scala 948:21]
  assign const12_io_enable_bits_taskID = bb_for_body3418_io_Out_1_bits_taskID; // @[extracted_function_reduction.scala 948:21]
  assign const12_io_Out_ready = binaryOp_inc68_io_RightIO_ready; // @[extracted_function_reduction.scala 1068:29]
  assign const13_clock = clock;
  assign const13_reset = reset;
  assign const13_io_enable_valid = bb_for_body3418_io_Out_2_valid; // @[extracted_function_reduction.scala 950:21]
  assign const13_io_enable_bits_taskID = bb_for_body3418_io_Out_2_bits_taskID; // @[extracted_function_reduction.scala 950:21]
  assign const13_io_Out_ready = icmp_exitcond69_io_RightIO_ready; // @[extracted_function_reduction.scala 1070:30]
endmodule

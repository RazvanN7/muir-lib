module LockingRRArbiter(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [15:0] io_in_0_bits_RouteID,
  input  [21:0] io_in_0_bits_address,
  input  [31:0] io_in_0_bits_data,
  input  [4:0]  io_in_0_bits_taskID,
  input  [7:0]  io_in_0_bits_Typ,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [15:0] io_in_1_bits_RouteID,
  input  [21:0] io_in_1_bits_address,
  input  [31:0] io_in_1_bits_data,
  input  [4:0]  io_in_1_bits_taskID,
  input  [7:0]  io_in_1_bits_Typ,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [21:0] io_out_bits_address,
  output [31:0] io_out_bits_data,
  output [4:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ,
  output        io_chosen
);
  wire  _T; // @[Decoupled.scala 40:37]
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Arbiter.scala 67:57]
  wire  _T_5; // @[Arbiter.scala 68:83]
  wire  _T_7; // @[Arbiter.scala 31:68]
  wire  _T_9; // @[Arbiter.scala 31:78]
  wire  _T_10; // @[Arbiter.scala 31:78]
  wire  _T_14; // @[Arbiter.scala 72:50]
  wire  _GEN_17; // @[Arbiter.scala 77:27]
  assign _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = 1'h1 > _T_1; // @[Arbiter.scala 67:57]
  assign _T_5 = io_in_1_valid & _T_3; // @[Arbiter.scala 68:83]
  assign _T_7 = _T_5 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_9 = _T_5 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_10 = _T_7 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_14 = _T_3 | _T_10; // @[Arbiter.scala 72:50]
  assign _GEN_17 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_9 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_14 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_RouteID = io_chosen ? io_in_1_bits_RouteID : io_in_0_bits_RouteID; // @[Arbiter.scala 42:15]
  assign io_out_bits_address = io_chosen ? io_in_1_bits_address : io_in_0_bits_address; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_out_bits_taskID = io_chosen ? io_in_1_bits_taskID : io_in_0_bits_taskID; // @[Arbiter.scala 42:15]
  assign io_out_bits_Typ = io_chosen ? io_in_1_bits_Typ : io_in_0_bits_Typ; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_5 | _GEN_17; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (_T) begin
      _T_1 <= io_chosen;
    end
  end
endmodule
module ArbiterTree(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [21:0] io_in_0_bits_address,
  input  [31:0] io_in_0_bits_data,
  input  [4:0]  io_in_0_bits_taskID,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [21:0] io_in_1_bits_address,
  input  [31:0] io_in_1_bits_data,
  input  [4:0]  io_in_1_bits_taskID,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [21:0] io_in_2_bits_address,
  input  [31:0] io_in_2_bits_data,
  input  [4:0]  io_in_2_bits_taskID,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [21:0] io_in_3_bits_address,
  input  [31:0] io_in_3_bits_data,
  input  [4:0]  io_in_3_bits_taskID,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [21:0] io_in_4_bits_address,
  input  [31:0] io_in_4_bits_data,
  input  [4:0]  io_in_4_bits_taskID,
  output        io_in_5_ready,
  input         io_in_5_valid,
  input  [21:0] io_in_5_bits_address,
  input  [31:0] io_in_5_bits_data,
  input  [4:0]  io_in_5_bits_taskID,
  output        io_in_6_ready,
  input         io_in_6_valid,
  input  [21:0] io_in_6_bits_address,
  input  [31:0] io_in_6_bits_data,
  input  [4:0]  io_in_6_bits_taskID,
  output        io_in_7_ready,
  input         io_in_7_valid,
  input  [21:0] io_in_7_bits_address,
  input  [31:0] io_in_7_bits_data,
  input  [4:0]  io_in_7_bits_taskID,
  output        io_in_8_ready,
  input         io_in_8_valid,
  input  [21:0] io_in_8_bits_address,
  input  [31:0] io_in_8_bits_data,
  input  [4:0]  io_in_8_bits_taskID,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [21:0] io_out_bits_address,
  output [31:0] io_out_bits_data,
  output [4:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ
);
  wire  LockingRRArbiter_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_1_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_1_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_1_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_1_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_1_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_1_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_1_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_1_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_1_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_1_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_1_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_1_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_1_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_1_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_1_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_2_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_2_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_2_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_2_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_2_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_2_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_2_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_2_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_2_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_2_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_2_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_2_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_2_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_2_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_2_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_3_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_3_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_3_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_3_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_3_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_3_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_3_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_3_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_3_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_3_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_3_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_3_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_3_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_3_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_3_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_4_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_4_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_4_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_4_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_4_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_4_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_4_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_4_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_4_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_4_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_4_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_4_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_4_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_4_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_4_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_5_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_5_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_5_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_5_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_5_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_5_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_5_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_5_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_5_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_5_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_5_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_5_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_5_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_5_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_5_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_6_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_6_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_6_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_6_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_6_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_6_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_6_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_6_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_6_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_6_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_6_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_6_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_6_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_6_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_6_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_7_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_7_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_7_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_7_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_7_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_7_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_7_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_7_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_7_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_7_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_7_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_7_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_7_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_7_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_7_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_8_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_8_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_8_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_8_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_8_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_8_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_8_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_8_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_8_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_8_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_8_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_8_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_8_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_8_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_8_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_9_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_9_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_9_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_9_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_9_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_9_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_9_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_9_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_9_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_9_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_9_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_9_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_9_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_9_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_9_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_10_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_10_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_10_io_in_0_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_10_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_10_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_10_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_10_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_10_io_in_1_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_10_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_10_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_10_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [21:0] LockingRRArbiter_10_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_10_io_out_bits_data; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_10_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_10_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_chosen; // @[ArbiterTree.scala 32:13]
  LockingRRArbiter LockingRRArbiter ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_clock),
    .io_in_0_ready(LockingRRArbiter_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_io_out_ready),
    .io_out_valid(LockingRRArbiter_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_1 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_1_clock),
    .io_in_0_ready(LockingRRArbiter_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_1_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_1_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_1_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_1_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_1_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_1_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_1_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_1_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_1_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_1_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_1_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_1_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_1_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_1_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_1_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_1_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_1_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_1_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_1_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_2 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_2_clock),
    .io_in_0_ready(LockingRRArbiter_2_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_2_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_2_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_2_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_2_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_2_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_2_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_2_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_2_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_2_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_2_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_2_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_2_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_2_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_2_io_out_ready),
    .io_out_valid(LockingRRArbiter_2_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_2_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_2_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_2_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_2_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_2_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_2_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_3 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_3_clock),
    .io_in_0_ready(LockingRRArbiter_3_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_3_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_3_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_3_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_3_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_3_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_3_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_3_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_3_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_3_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_3_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_3_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_3_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_3_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_3_io_out_ready),
    .io_out_valid(LockingRRArbiter_3_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_3_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_3_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_3_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_3_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_3_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_3_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_4 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_4_clock),
    .io_in_0_ready(LockingRRArbiter_4_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_4_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_4_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_4_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_4_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_4_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_4_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_4_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_4_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_4_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_4_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_4_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_4_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_4_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_4_io_out_ready),
    .io_out_valid(LockingRRArbiter_4_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_4_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_4_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_4_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_4_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_4_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_4_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_5 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_5_clock),
    .io_in_0_ready(LockingRRArbiter_5_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_5_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_5_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_5_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_5_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_5_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_5_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_5_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_5_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_5_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_5_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_5_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_5_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_5_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_5_io_out_ready),
    .io_out_valid(LockingRRArbiter_5_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_5_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_5_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_5_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_5_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_5_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_5_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_6 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_6_clock),
    .io_in_0_ready(LockingRRArbiter_6_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_6_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_6_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_6_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_6_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_6_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_6_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_6_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_6_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_6_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_6_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_6_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_6_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_6_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_6_io_out_ready),
    .io_out_valid(LockingRRArbiter_6_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_6_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_6_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_6_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_6_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_6_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_6_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_7 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_7_clock),
    .io_in_0_ready(LockingRRArbiter_7_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_7_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_7_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_7_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_7_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_7_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_7_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_7_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_7_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_7_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_7_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_7_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_7_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_7_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_7_io_out_ready),
    .io_out_valid(LockingRRArbiter_7_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_7_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_7_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_7_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_7_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_7_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_7_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_8 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_8_clock),
    .io_in_0_ready(LockingRRArbiter_8_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_8_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_8_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_8_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_8_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_8_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_8_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_8_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_8_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_8_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_8_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_8_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_8_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_8_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_8_io_out_ready),
    .io_out_valid(LockingRRArbiter_8_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_8_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_8_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_8_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_8_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_8_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_8_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_9 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_9_clock),
    .io_in_0_ready(LockingRRArbiter_9_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_9_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_9_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_9_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_9_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_9_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_9_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_9_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_9_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_9_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_9_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_9_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_9_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_9_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_9_io_out_ready),
    .io_out_valid(LockingRRArbiter_9_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_9_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_9_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_9_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_9_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_9_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_9_io_chosen)
  );
  LockingRRArbiter LockingRRArbiter_10 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_10_clock),
    .io_in_0_ready(LockingRRArbiter_10_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_10_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_10_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_10_io_in_0_bits_address),
    .io_in_0_bits_data(LockingRRArbiter_10_io_in_0_bits_data),
    .io_in_0_bits_taskID(LockingRRArbiter_10_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_10_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_10_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_10_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_10_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_10_io_in_1_bits_address),
    .io_in_1_bits_data(LockingRRArbiter_10_io_in_1_bits_data),
    .io_in_1_bits_taskID(LockingRRArbiter_10_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_10_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_10_io_out_ready),
    .io_out_valid(LockingRRArbiter_10_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_10_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_10_io_out_bits_address),
    .io_out_bits_data(LockingRRArbiter_10_io_out_bits_data),
    .io_out_bits_taskID(LockingRRArbiter_10_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_10_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_10_io_chosen)
  );
  assign io_in_0_ready = LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_1_ready = LockingRRArbiter_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_2_ready = LockingRRArbiter_1_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_3_ready = LockingRRArbiter_1_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_4_ready = LockingRRArbiter_2_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_5_ready = LockingRRArbiter_2_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_6_ready = LockingRRArbiter_3_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_7_ready = LockingRRArbiter_3_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_8_ready = LockingRRArbiter_4_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_out_valid = LockingRRArbiter_10_io_out_valid; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_RouteID = LockingRRArbiter_10_io_out_bits_RouteID; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_address = LockingRRArbiter_10_io_out_bits_address; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_data = LockingRRArbiter_10_io_out_bits_data; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_taskID = LockingRRArbiter_10_io_out_bits_taskID; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_Typ = LockingRRArbiter_10_io_out_bits_Typ; // @[ArbiterTree.scala 65:12]
  assign LockingRRArbiter_clock = clock;
  assign LockingRRArbiter_io_in_0_valid = io_in_0_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_RouteID = 16'h0; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_address = io_in_0_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_data = io_in_0_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_taskID = io_in_0_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_valid = io_in_1_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_RouteID = 16'h1; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_address = io_in_1_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_data = io_in_1_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_taskID = io_in_1_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_out_ready = LockingRRArbiter_5_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_1_clock = clock;
  assign LockingRRArbiter_1_io_in_0_valid = io_in_2_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_RouteID = 16'h2; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_address = io_in_2_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_data = io_in_2_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_taskID = io_in_2_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_valid = io_in_3_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_bits_RouteID = 16'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_bits_address = io_in_3_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_bits_data = io_in_3_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_bits_taskID = io_in_3_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_out_ready = LockingRRArbiter_5_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_clock = clock;
  assign LockingRRArbiter_2_io_in_0_valid = io_in_4_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_0_bits_RouteID = 16'h4; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_0_bits_address = io_in_4_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_0_bits_data = io_in_4_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_0_bits_taskID = io_in_4_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_valid = io_in_5_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_bits_RouteID = 16'h5; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_bits_address = io_in_5_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_bits_data = io_in_5_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_bits_taskID = io_in_5_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_out_ready = LockingRRArbiter_6_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_3_clock = clock;
  assign LockingRRArbiter_3_io_in_0_valid = io_in_6_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_0_bits_RouteID = 16'h6; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_0_bits_address = io_in_6_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_0_bits_data = io_in_6_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_0_bits_taskID = io_in_6_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_valid = io_in_7_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_bits_RouteID = 16'h7; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_bits_address = io_in_7_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_bits_data = io_in_7_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_bits_taskID = io_in_7_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_out_ready = LockingRRArbiter_6_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_4_clock = clock;
  assign LockingRRArbiter_4_io_in_0_valid = io_in_8_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_0_bits_RouteID = 16'h8; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_0_bits_address = io_in_8_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_0_bits_data = io_in_8_bits_data; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_0_bits_taskID = io_in_8_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_1_valid = 1'h0; // @[ArbiterTree.scala 52:67]
  assign LockingRRArbiter_4_io_in_1_bits_RouteID = 16'h0;
  assign LockingRRArbiter_4_io_in_1_bits_address = 22'h0;
  assign LockingRRArbiter_4_io_in_1_bits_data = 32'h0;
  assign LockingRRArbiter_4_io_in_1_bits_taskID = 5'h0;
  assign LockingRRArbiter_4_io_in_1_bits_Typ = 8'h0;
  assign LockingRRArbiter_4_io_out_ready = LockingRRArbiter_7_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_clock = clock;
  assign LockingRRArbiter_5_io_in_0_valid = LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_0_bits_RouteID = LockingRRArbiter_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_0_bits_address = LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_0_bits_data = LockingRRArbiter_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_0_bits_taskID = LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_0_bits_Typ = LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_1_valid = LockingRRArbiter_1_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_1_bits_RouteID = LockingRRArbiter_1_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_1_bits_address = LockingRRArbiter_1_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_1_bits_data = LockingRRArbiter_1_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_1_bits_taskID = LockingRRArbiter_1_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_in_1_bits_Typ = LockingRRArbiter_1_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_io_out_ready = LockingRRArbiter_8_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_clock = clock;
  assign LockingRRArbiter_6_io_in_0_valid = LockingRRArbiter_2_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_0_bits_RouteID = LockingRRArbiter_2_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_0_bits_address = LockingRRArbiter_2_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_0_bits_data = LockingRRArbiter_2_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_0_bits_taskID = LockingRRArbiter_2_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_0_bits_Typ = LockingRRArbiter_2_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_1_valid = LockingRRArbiter_3_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_1_bits_RouteID = LockingRRArbiter_3_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_1_bits_address = LockingRRArbiter_3_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_1_bits_data = LockingRRArbiter_3_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_1_bits_taskID = LockingRRArbiter_3_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_in_1_bits_Typ = LockingRRArbiter_3_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_io_out_ready = LockingRRArbiter_8_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_7_clock = clock;
  assign LockingRRArbiter_7_io_in_0_valid = LockingRRArbiter_4_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_7_io_in_0_bits_RouteID = LockingRRArbiter_4_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_7_io_in_0_bits_address = LockingRRArbiter_4_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_7_io_in_0_bits_data = LockingRRArbiter_4_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_7_io_in_0_bits_taskID = LockingRRArbiter_4_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_7_io_in_0_bits_Typ = LockingRRArbiter_4_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_7_io_in_1_valid = 1'h0; // @[ArbiterTree.scala 39:67]
  assign LockingRRArbiter_7_io_in_1_bits_RouteID = 16'h0;
  assign LockingRRArbiter_7_io_in_1_bits_address = 22'h0;
  assign LockingRRArbiter_7_io_in_1_bits_data = 32'h0;
  assign LockingRRArbiter_7_io_in_1_bits_taskID = 5'h0;
  assign LockingRRArbiter_7_io_in_1_bits_Typ = 8'h0;
  assign LockingRRArbiter_7_io_out_ready = LockingRRArbiter_9_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_clock = clock;
  assign LockingRRArbiter_8_io_in_0_valid = LockingRRArbiter_5_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_0_bits_RouteID = LockingRRArbiter_5_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_0_bits_address = LockingRRArbiter_5_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_0_bits_data = LockingRRArbiter_5_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_0_bits_taskID = LockingRRArbiter_5_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_0_bits_Typ = LockingRRArbiter_5_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_1_valid = LockingRRArbiter_6_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_1_bits_RouteID = LockingRRArbiter_6_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_1_bits_address = LockingRRArbiter_6_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_1_bits_data = LockingRRArbiter_6_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_1_bits_taskID = LockingRRArbiter_6_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_in_1_bits_Typ = LockingRRArbiter_6_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_io_out_ready = LockingRRArbiter_10_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_9_clock = clock;
  assign LockingRRArbiter_9_io_in_0_valid = LockingRRArbiter_7_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_9_io_in_0_bits_RouteID = LockingRRArbiter_7_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_9_io_in_0_bits_address = LockingRRArbiter_7_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_9_io_in_0_bits_data = LockingRRArbiter_7_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_9_io_in_0_bits_taskID = LockingRRArbiter_7_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_9_io_in_0_bits_Typ = LockingRRArbiter_7_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_9_io_in_1_valid = 1'h0; // @[ArbiterTree.scala 39:67]
  assign LockingRRArbiter_9_io_in_1_bits_RouteID = 16'h0;
  assign LockingRRArbiter_9_io_in_1_bits_address = 22'h0;
  assign LockingRRArbiter_9_io_in_1_bits_data = 32'h0;
  assign LockingRRArbiter_9_io_in_1_bits_taskID = 5'h0;
  assign LockingRRArbiter_9_io_in_1_bits_Typ = 8'h0;
  assign LockingRRArbiter_9_io_out_ready = LockingRRArbiter_10_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_clock = clock;
  assign LockingRRArbiter_10_io_in_0_valid = LockingRRArbiter_8_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_0_bits_RouteID = LockingRRArbiter_8_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_0_bits_address = LockingRRArbiter_8_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_0_bits_data = LockingRRArbiter_8_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_0_bits_taskID = LockingRRArbiter_8_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_0_bits_Typ = LockingRRArbiter_8_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_valid = LockingRRArbiter_9_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_bits_RouteID = LockingRRArbiter_9_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_bits_address = LockingRRArbiter_9_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_bits_data = LockingRRArbiter_9_io_out_bits_data; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_bits_taskID = LockingRRArbiter_9_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_bits_Typ = LockingRRArbiter_9_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_out_ready = io_out_ready; // @[ArbiterTree.scala 65:12]
endmodule
module Arbiter(
  output  io_in_0_ready,
  input   io_in_0_valid,
  output  io_in_1_ready,
  input   io_in_1_valid,
  input   io_out_ready,
  output  io_out_valid
);
  wire  _T; // @[Arbiter.scala 31:78]
  wire  _T_3; // @[Arbiter.scala 135:19]
  assign _T = io_in_0_valid == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_3 = _T == 1'h0; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = _T & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_3 | io_in_1_valid; // @[Arbiter.scala 135:16]
endmodule
module Arbiter_1(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [31:0] io_in_0_bits_data,
  input  [3:0]  io_in_0_bits_mask,
  input  [7:0]  io_in_0_bits_tag,
  input  [4:0]  io_in_0_bits_taskID,
  input         io_in_0_bits_iswrite,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [31:0] io_in_1_bits_data,
  input  [3:0]  io_in_1_bits_mask,
  input  [7:0]  io_in_1_bits_tag,
  input  [4:0]  io_in_1_bits_taskID,
  input         io_in_1_bits_iswrite,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [31:0] io_out_bits_data,
  output [3:0]  io_out_bits_mask,
  output [7:0]  io_out_bits_tag,
  output [4:0]  io_out_bits_taskID,
  output        io_out_bits_iswrite
);
  wire  _T; // @[Arbiter.scala 31:78]
  wire  _T_3; // @[Arbiter.scala 135:19]
  assign _T = io_in_0_valid == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_3 = _T == 1'h0; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = _T & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_3 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : io_in_1_bits_data; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_mask = io_in_0_valid ? io_in_0_bits_mask : io_in_1_bits_mask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_tag = io_in_0_valid ? io_in_0_bits_tag : io_in_1_bits_tag; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_taskID = io_in_0_valid ? io_in_0_bits_taskID : io_in_1_bits_taskID; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_iswrite = io_in_0_valid ? io_in_0_bits_iswrite : io_in_1_bits_iswrite; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Demux(
  input         io_en,
  input  [31:0] io_input_data,
  input  [7:0]  io_input_tag,
  input         io_sel,
  output        io_outputs_0_valid,
  output [31:0] io_outputs_0_data,
  output [7:0]  io_outputs_0_tag,
  output        io_outputs_1_valid,
  output [31:0] io_outputs_1_data,
  output [7:0]  io_outputs_1_tag
);
  wire  _GEN_0; // @[Muxes.scala 29:25]
  assign _GEN_0 = 1'h0 == io_sel; // @[Muxes.scala 29:25]
  assign io_outputs_0_valid = io_en & _GEN_0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_0_data = io_input_data; // @[Muxes.scala 23:19]
  assign io_outputs_0_tag = io_input_tag; // @[Muxes.scala 23:19]
  assign io_outputs_1_valid = io_en & io_sel; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_1_data = io_input_data; // @[Muxes.scala 23:19]
  assign io_outputs_1_tag = io_input_tag; // @[Muxes.scala 23:19]
endmodule
module RRArbiter(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [15:0] io_in_0_bits_RouteID,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [15:0] io_in_1_bits_RouteID,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output        io_chosen
);
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Arbiter.scala 67:57]
  wire  _T_5; // @[Arbiter.scala 68:83]
  wire  _T_7; // @[Arbiter.scala 31:68]
  wire  _T_10; // @[Arbiter.scala 31:78]
  wire  _GEN_11; // @[Arbiter.scala 77:27]
  assign _T_3 = 1'h1 > _T_1; // @[Arbiter.scala 67:57]
  assign _T_5 = io_in_1_valid & _T_3; // @[Arbiter.scala 68:83]
  assign _T_7 = _T_5 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_10 = _T_7 == 1'h0; // @[Arbiter.scala 31:78]
  assign _GEN_11 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_5 == 1'h0; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_3 | _T_10; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_RouteID = io_chosen ? io_in_1_bits_RouteID : io_in_0_bits_RouteID; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_5 | _GEN_11; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_out_valid) begin
      _T_1 <= io_chosen;
    end
  end
endmodule
module Demux_1(
  input         io_en,
  input  [15:0] io_input_RouteID,
  input         io_sel,
  output        io_outputs_0_valid,
  output [15:0] io_outputs_0_RouteID,
  output        io_outputs_1_valid,
  output [15:0] io_outputs_1_RouteID
);
  wire  _GEN_0; // @[Muxes.scala 29:25]
  assign _GEN_0 = 1'h0 == io_sel; // @[Muxes.scala 29:25]
  assign io_outputs_0_valid = io_en & _GEN_0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_0_RouteID = io_input_RouteID; // @[Muxes.scala 23:19]
  assign io_outputs_1_valid = io_en & io_sel; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_1_RouteID = io_input_RouteID; // @[Muxes.scala 23:19]
endmodule
module DeMuxTree(
  input         clock,
  input         reset,
  output        io_outputs_0_valid,
  output        io_outputs_1_valid,
  output        io_outputs_2_valid,
  output        io_outputs_3_valid,
  output        io_outputs_4_valid,
  output        io_outputs_5_valid,
  output        io_outputs_6_valid,
  output        io_outputs_7_valid,
  output        io_outputs_8_valid,
  input  [15:0] io_input_RouteID,
  input         io_enable
);
  wire  Demux_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_1_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_1_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_1_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_1_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_1_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_1_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_1_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_2_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_2_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_2_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_2_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_2_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_2_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_2_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_3_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_3_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_3_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_3_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_3_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_3_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_3_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_4_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_4_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_4_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_4_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_4_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_4_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_4_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_5_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_5_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_5_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_5_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_5_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_5_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_5_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_6_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_6_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_6_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_6_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_6_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_6_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_6_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_7_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_7_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_7_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_7_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_7_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_7_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_7_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_8_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_8_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_8_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_8_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_8_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_8_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_8_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_9_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_9_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_9_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_9_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_9_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_9_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_9_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_10_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_10_io_input_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_10_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_10_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_10_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire  Demux_10_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_10_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  reg [15:0] _T_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_1;
  reg [15:0] _T_3_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_2;
  reg  _T_4; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_3;
  reg [15:0] _T_6_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_4;
  reg  _T_7; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_5;
  reg [15:0] _T_9_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_6;
  reg  _T_10; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_7;
  reg [15:0] _T_12_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_8;
  reg  _T_13; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_9;
  reg [15:0] _T_15_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_10;
  reg  _T_16; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_11;
  reg [15:0] _T_18_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_12;
  reg  _T_19; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_13;
  reg [15:0] _T_21_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_14;
  reg  _T_22; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_15;
  reg [15:0] _T_24_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_16;
  reg  _T_25; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_17;
  reg [15:0] _T_27_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_18;
  reg  _T_28; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_19;
  Demux_1 Demux ( // @[Muxes.scala 91:13]
    .io_en(Demux_io_en),
    .io_input_RouteID(Demux_io_input_RouteID),
    .io_sel(Demux_io_sel),
    .io_outputs_0_valid(Demux_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_io_outputs_1_RouteID)
  );
  Demux_1 Demux_1 ( // @[Muxes.scala 91:13]
    .io_en(Demux_1_io_en),
    .io_input_RouteID(Demux_1_io_input_RouteID),
    .io_sel(Demux_1_io_sel),
    .io_outputs_0_valid(Demux_1_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_1_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_1_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_1_io_outputs_1_RouteID)
  );
  Demux_1 Demux_2 ( // @[Muxes.scala 91:13]
    .io_en(Demux_2_io_en),
    .io_input_RouteID(Demux_2_io_input_RouteID),
    .io_sel(Demux_2_io_sel),
    .io_outputs_0_valid(Demux_2_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_2_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_2_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_2_io_outputs_1_RouteID)
  );
  Demux_1 Demux_3 ( // @[Muxes.scala 91:13]
    .io_en(Demux_3_io_en),
    .io_input_RouteID(Demux_3_io_input_RouteID),
    .io_sel(Demux_3_io_sel),
    .io_outputs_0_valid(Demux_3_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_3_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_3_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_3_io_outputs_1_RouteID)
  );
  Demux_1 Demux_4 ( // @[Muxes.scala 91:13]
    .io_en(Demux_4_io_en),
    .io_input_RouteID(Demux_4_io_input_RouteID),
    .io_sel(Demux_4_io_sel),
    .io_outputs_0_valid(Demux_4_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_4_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_4_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_4_io_outputs_1_RouteID)
  );
  Demux_1 Demux_5 ( // @[Muxes.scala 91:13]
    .io_en(Demux_5_io_en),
    .io_input_RouteID(Demux_5_io_input_RouteID),
    .io_sel(Demux_5_io_sel),
    .io_outputs_0_valid(Demux_5_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_5_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_5_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_5_io_outputs_1_RouteID)
  );
  Demux_1 Demux_6 ( // @[Muxes.scala 91:13]
    .io_en(Demux_6_io_en),
    .io_input_RouteID(Demux_6_io_input_RouteID),
    .io_sel(Demux_6_io_sel),
    .io_outputs_0_valid(Demux_6_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_6_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_6_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_6_io_outputs_1_RouteID)
  );
  Demux_1 Demux_7 ( // @[Muxes.scala 91:13]
    .io_en(Demux_7_io_en),
    .io_input_RouteID(Demux_7_io_input_RouteID),
    .io_sel(Demux_7_io_sel),
    .io_outputs_0_valid(Demux_7_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_7_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_7_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_7_io_outputs_1_RouteID)
  );
  Demux_1 Demux_8 ( // @[Muxes.scala 91:13]
    .io_en(Demux_8_io_en),
    .io_input_RouteID(Demux_8_io_input_RouteID),
    .io_sel(Demux_8_io_sel),
    .io_outputs_0_valid(Demux_8_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_8_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_8_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_8_io_outputs_1_RouteID)
  );
  Demux_1 Demux_9 ( // @[Muxes.scala 91:13]
    .io_en(Demux_9_io_en),
    .io_input_RouteID(Demux_9_io_input_RouteID),
    .io_sel(Demux_9_io_sel),
    .io_outputs_0_valid(Demux_9_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_9_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_9_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_9_io_outputs_1_RouteID)
  );
  Demux_1 Demux_10 ( // @[Muxes.scala 91:13]
    .io_en(Demux_10_io_en),
    .io_input_RouteID(Demux_10_io_input_RouteID),
    .io_sel(Demux_10_io_sel),
    .io_outputs_0_valid(Demux_10_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_10_io_outputs_0_RouteID),
    .io_outputs_1_valid(Demux_10_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_10_io_outputs_1_RouteID)
  );
  assign io_outputs_0_valid = Demux_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_1_valid = Demux_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_2_valid = Demux_1_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_3_valid = Demux_1_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_4_valid = Demux_2_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_5_valid = Demux_2_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_6_valid = Demux_3_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_7_valid = Demux_3_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_8_valid = Demux_4_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign Demux_io_en = _T_1; // @[Muxes.scala 105:20]
  assign Demux_io_input_RouteID = _T_RouteID; // @[Muxes.scala 104:23]
  assign Demux_io_sel = _T_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_1_io_en = _T_4; // @[Muxes.scala 105:20]
  assign Demux_1_io_input_RouteID = _T_3_RouteID; // @[Muxes.scala 104:23]
  assign Demux_1_io_sel = _T_3_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_2_io_en = _T_7; // @[Muxes.scala 105:20]
  assign Demux_2_io_input_RouteID = _T_6_RouteID; // @[Muxes.scala 104:23]
  assign Demux_2_io_sel = _T_6_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_3_io_en = _T_10; // @[Muxes.scala 105:20]
  assign Demux_3_io_input_RouteID = _T_9_RouteID; // @[Muxes.scala 104:23]
  assign Demux_3_io_sel = _T_9_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_4_io_en = _T_13; // @[Muxes.scala 105:20]
  assign Demux_4_io_input_RouteID = _T_12_RouteID; // @[Muxes.scala 104:23]
  assign Demux_4_io_sel = _T_12_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_5_io_en = _T_16; // @[Muxes.scala 105:20]
  assign Demux_5_io_input_RouteID = _T_15_RouteID; // @[Muxes.scala 104:23]
  assign Demux_5_io_sel = _T_15_RouteID[1]; // @[Muxes.scala 106:21]
  assign Demux_6_io_en = _T_19; // @[Muxes.scala 105:20]
  assign Demux_6_io_input_RouteID = _T_18_RouteID; // @[Muxes.scala 104:23]
  assign Demux_6_io_sel = _T_18_RouteID[1]; // @[Muxes.scala 106:21]
  assign Demux_7_io_en = _T_22; // @[Muxes.scala 105:20]
  assign Demux_7_io_input_RouteID = _T_21_RouteID; // @[Muxes.scala 104:23]
  assign Demux_7_io_sel = _T_21_RouteID[1]; // @[Muxes.scala 106:21]
  assign Demux_8_io_en = _T_25; // @[Muxes.scala 105:20]
  assign Demux_8_io_input_RouteID = _T_24_RouteID; // @[Muxes.scala 104:23]
  assign Demux_8_io_sel = _T_24_RouteID[2]; // @[Muxes.scala 106:21]
  assign Demux_9_io_en = _T_28; // @[Muxes.scala 105:20]
  assign Demux_9_io_input_RouteID = _T_27_RouteID; // @[Muxes.scala 104:23]
  assign Demux_9_io_sel = _T_27_RouteID[2]; // @[Muxes.scala 106:21]
  assign Demux_10_io_en = io_enable; // @[Muxes.scala 135:14]
  assign Demux_10_io_input_RouteID = io_input_RouteID; // @[Muxes.scala 134:17]
  assign Demux_10_io_sel = io_input_RouteID[3]; // @[Muxes.scala 136:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_RouteID = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_3_RouteID = _RAND_2[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_4 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_6_RouteID = _RAND_4[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_7 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_9_RouteID = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_10 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_12_RouteID = _RAND_8[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_13 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_15_RouteID = _RAND_10[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_16 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_18_RouteID = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_19 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_21_RouteID = _RAND_14[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_22 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_24_RouteID = _RAND_16[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_25 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_27_RouteID = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_28 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    _T_RouteID <= Demux_5_io_outputs_0_RouteID;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= Demux_5_io_outputs_0_valid;
    end
    _T_3_RouteID <= Demux_5_io_outputs_1_RouteID;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= Demux_5_io_outputs_1_valid;
    end
    _T_6_RouteID <= Demux_6_io_outputs_0_RouteID;
    if (reset) begin
      _T_7 <= 1'h0;
    end else begin
      _T_7 <= Demux_6_io_outputs_0_valid;
    end
    _T_9_RouteID <= Demux_6_io_outputs_1_RouteID;
    if (reset) begin
      _T_10 <= 1'h0;
    end else begin
      _T_10 <= Demux_6_io_outputs_1_valid;
    end
    _T_12_RouteID <= Demux_7_io_outputs_0_RouteID;
    if (reset) begin
      _T_13 <= 1'h0;
    end else begin
      _T_13 <= Demux_7_io_outputs_0_valid;
    end
    _T_15_RouteID <= Demux_8_io_outputs_0_RouteID;
    if (reset) begin
      _T_16 <= 1'h0;
    end else begin
      _T_16 <= Demux_8_io_outputs_0_valid;
    end
    _T_18_RouteID <= Demux_8_io_outputs_1_RouteID;
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      _T_19 <= Demux_8_io_outputs_1_valid;
    end
    _T_21_RouteID <= Demux_9_io_outputs_0_RouteID;
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      _T_22 <= Demux_9_io_outputs_0_valid;
    end
    _T_24_RouteID <= Demux_10_io_outputs_0_RouteID;
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      _T_25 <= Demux_10_io_outputs_0_valid;
    end
    _T_27_RouteID <= Demux_10_io_outputs_1_RouteID;
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      _T_28 <= Demux_10_io_outputs_1_valid;
    end
  end
endmodule
module WriteTableEntry(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [15:0] io_NodeReq_bits_RouteID,
  input  [21:0] io_NodeReq_bits_address,
  input  [31:0] io_NodeReq_bits_data,
  input  [4:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output        io_free
);
  reg [15:0] request_R_RouteID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_0;
  reg [4:0] request_R_taskID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_1;
  reg [7:0] sendbytemask; // @[WriteMemoryController.scala 61:29]
  reg [31:0] _RAND_2;
  reg [31:0] ReqAddress; // @[WriteMemoryController.scala 65:27]
  reg [31:0] _RAND_3;
  reg  ptr; // @[WriteMemoryController.scala 70:27]
  reg [31:0] _RAND_4;
  reg [31:0] linebuffer_0; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_5;
  reg [31:0] linebuffer_1; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_6;
  reg [1:0] state; // @[WriteMemoryController.scala 76:68]
  reg [31:0] _RAND_7;
  wire  _T_4; // @[WriteMemoryController.scala 89:21]
  wire [2:0] _T_5; // @[Cat.scala 29:58]
  wire [31:0] _GEN_29; // @[WriteMemoryController.scala 100:37]
  reg  isWrite; // @[WriteMemoryController.scala 108:24]
  reg [31:0] _RAND_8;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire [19:0] _T_10; // @[WriteMemoryController.scala 121:44]
  wire [21:0] _T_11; // @[WriteMemoryController.scala 121:69]
  wire  _T_12; // @[helpers.scala 27:24]
  wire  _T_13; // @[helpers.scala 27:47]
  wire  _T_14; // @[helpers.scala 27:40]
  wire  _T_16; // @[helpers.scala 28:15]
  wire  _T_17; // @[helpers.scala 28:38]
  wire  _T_18; // @[helpers.scala 28:31]
  wire  _T_20; // @[helpers.scala 29:17]
  wire  _T_21; // @[helpers.scala 29:40]
  wire  _T_22; // @[helpers.scala 29:33]
  wire [1:0] _T_28; // @[helpers.scala 39:32]
  wire [4:0] _T_29; // @[Cat.scala 29:58]
  wire [7:0] _T_43; // @[helpers.scala 50:12]
  wire [7:0] _T_44; // @[helpers.scala 49:10]
  wire [7:0] _T_45; // @[helpers.scala 48:19]
  wire [10:0] _GEN_31; // @[helpers.scala 20:26]
  wire [10:0] _T_47; // @[helpers.scala 20:26]
  wire [62:0] _GEN_32; // @[WriteMemoryController.scala 127:41]
  wire [62:0] _T_50; // @[WriteMemoryController.scala 127:41]
  wire [63:0] _T_52;
  wire [31:0] _T_53; // @[WriteMemoryController.scala 127:121]
  wire [31:0] _T_54; // @[WriteMemoryController.scala 127:121]
  wire [10:0] _GEN_10; // @[WriteMemoryController.scala 117:28]
  wire  _T_55; // @[WriteMemoryController.scala 139:15]
  wire  _T_56; // @[WriteMemoryController.scala 139:47]
  wire  _T_57; // @[WriteMemoryController.scala 139:30]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire [3:0] _T_59; // @[WriteMemoryController.scala 144:36]
  wire  _T_61; // @[WriteMemoryController.scala 146:18]
  wire [10:0] _GEN_14; // @[WriteMemoryController.scala 142:29]
  wire [10:0] _GEN_18; // @[WriteMemoryController.scala 139:76]
  wire  _T_62; // @[WriteMemoryController.scala 156:15]
  wire  _T_64; // @[WriteMemoryController.scala 156:32]
  wire  _T_65; // @[WriteMemoryController.scala 158:27]
  wire  _T_68; // @[Decoupled.scala 40:37]
  assign _T_4 = state == 2'h3; // @[WriteMemoryController.scala 89:21]
  assign _T_5 = {ptr,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_29 = {{29'd0}, _T_5}; // @[WriteMemoryController.scala 100:37]
  assign _T_9 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_NodeReq_bits_address[21:2]; // @[WriteMemoryController.scala 121:44]
  assign _T_11 = {_T_10, 2'h0}; // @[WriteMemoryController.scala 121:69]
  assign _T_12 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_13 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_14 = _T_12 | _T_13; // @[helpers.scala 27:40]
  assign _T_16 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_17 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_18 = _T_16 | _T_17; // @[helpers.scala 28:31]
  assign _T_20 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_21 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_22 = _T_20 | _T_21; // @[helpers.scala 29:33]
  assign _T_28 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_29 = {_T_28,3'h0}; // @[Cat.scala 29:58]
  assign _T_43 = _T_22 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_44 = _T_18 ? 8'h1 : _T_43; // @[helpers.scala 49:10]
  assign _T_45 = _T_14 ? 8'h3 : _T_44; // @[helpers.scala 48:19]
  assign _GEN_31 = {{3'd0}, _T_45}; // @[helpers.scala 20:26]
  assign _T_47 = _GEN_31 << _T_28; // @[helpers.scala 20:26]
  assign _GEN_32 = {{31'd0}, io_NodeReq_bits_data}; // @[WriteMemoryController.scala 127:41]
  assign _T_50 = _GEN_32 << _T_29; // @[WriteMemoryController.scala 127:41]
  assign _T_52 = {{1'd0}, _T_50};
  assign _T_53 = _T_52[31:0]; // @[WriteMemoryController.scala 127:121]
  assign _T_54 = _T_52[63:32]; // @[WriteMemoryController.scala 127:121]
  assign _GEN_10 = _T_9 ? _T_47 : {{3'd0}, sendbytemask}; // @[WriteMemoryController.scala 117:28]
  assign _T_55 = state == 2'h1; // @[WriteMemoryController.scala 139:15]
  assign _T_56 = sendbytemask != 8'h0; // @[WriteMemoryController.scala 139:47]
  assign _T_57 = _T_55 & _T_56; // @[WriteMemoryController.scala 139:30]
  assign _T_58 = io_MemReq_ready & io_MemReq_valid; // @[Decoupled.scala 40:37]
  assign _T_59 = sendbytemask[7:4]; // @[WriteMemoryController.scala 144:36]
  assign _T_61 = ptr + 1'h1; // @[WriteMemoryController.scala 146:18]
  assign _GEN_14 = _T_58 ? {{7'd0}, _T_59} : _GEN_10; // @[WriteMemoryController.scala 142:29]
  assign _GEN_18 = _T_57 ? _GEN_14 : _GEN_10; // @[WriteMemoryController.scala 139:76]
  assign _T_62 = state == 2'h2; // @[WriteMemoryController.scala 156:15]
  assign _T_64 = _T_62 & io_MemResp_valid; // @[WriteMemoryController.scala 156:32]
  assign _T_65 = sendbytemask == 8'h0; // @[WriteMemoryController.scala 158:27]
  assign _T_68 = io_output_ready & io_output_valid; // @[Decoupled.scala 40:37]
  assign io_NodeReq_ready = state == 2'h0; // @[WriteMemoryController.scala 87:20]
  assign io_MemReq_valid = _T_55 & _T_56; // @[WriteMemoryController.scala 99:19 WriteMemoryController.scala 140:21]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_29; // @[WriteMemoryController.scala 100:23]
  assign io_MemReq_bits_data = ptr ? linebuffer_1 : linebuffer_0; // @[WriteMemoryController.scala 102:23]
  assign io_MemReq_bits_mask = sendbytemask[3:0]; // @[WriteMemoryController.scala 103:23]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[WriteMemoryController.scala 110:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[WriteMemoryController.scala 109:26]
  assign io_output_valid = state == 2'h3; // @[WriteMemoryController.scala 95:19 WriteMemoryController.scala 168:21]
  assign io_output_bits_RouteID = request_R_RouteID; // @[WriteMemoryController.scala 98:26]
  assign io_free = state == 2'h0; // @[WriteMemoryController.scala 85:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  request_R_RouteID = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  sendbytemask = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ReqAddress = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ptr = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  linebuffer_0 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  linebuffer_1 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  isWrite = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_9) begin
        request_R_RouteID <= io_NodeReq_bits_RouteID;
      end
    end
    if (reset) begin
      request_R_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_18[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_9) begin
        ReqAddress <= {{10'd0}, _T_11};
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (_T_4) begin
        ptr <= 1'h0;
      end else begin
        if (_T_57) begin
          if (_T_58) begin
            ptr <= _T_61;
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (_T_9) begin
        linebuffer_0 <= _T_53;
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (_T_9) begin
        linebuffer_1 <= _T_54;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_4) begin
        if (_T_68) begin
          state <= 2'h0;
        end else begin
          if (_T_64) begin
            if (_T_65) begin
              state <= 2'h3;
            end else begin
              state <= 2'h1;
            end
          end else begin
            if (_T_57) begin
              if (_T_58) begin
                state <= 2'h2;
              end else begin
                if (_T_9) begin
                  state <= 2'h1;
                end
              end
            end else begin
              if (_T_9) begin
                state <= 2'h1;
              end
            end
          end
        end
      end else begin
        if (_T_64) begin
          if (_T_65) begin
            state <= 2'h3;
          end else begin
            state <= 2'h1;
          end
        end else begin
          if (_T_57) begin
            if (_T_58) begin
              state <= 2'h2;
            end else begin
              if (_T_9) begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_9) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      isWrite <= 1'h0;
    end else begin
      isWrite <= 1'h1;
    end
  end
endmodule
module WriteTableEntry_1(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [15:0] io_NodeReq_bits_RouteID,
  input  [21:0] io_NodeReq_bits_address,
  input  [31:0] io_NodeReq_bits_data,
  input  [4:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output        io_free
);
  reg  ID; // @[WriteMemoryController.scala 53:32]
  reg [31:0] _RAND_0;
  reg [15:0] request_R_RouteID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_1;
  reg [4:0] request_R_taskID; // @[WriteMemoryController.scala 54:32]
  reg [31:0] _RAND_2;
  reg [7:0] sendbytemask; // @[WriteMemoryController.scala 61:29]
  reg [31:0] _RAND_3;
  reg [31:0] ReqAddress; // @[WriteMemoryController.scala 65:27]
  reg [31:0] _RAND_4;
  reg  ptr; // @[WriteMemoryController.scala 70:27]
  reg [31:0] _RAND_5;
  reg [31:0] linebuffer_0; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_6;
  reg [31:0] linebuffer_1; // @[WriteMemoryController.scala 71:27]
  reg [31:0] _RAND_7;
  reg [1:0] state; // @[WriteMemoryController.scala 76:68]
  reg [31:0] _RAND_8;
  wire  _T_4; // @[WriteMemoryController.scala 89:21]
  wire [2:0] _T_5; // @[Cat.scala 29:58]
  wire [31:0] _GEN_29; // @[WriteMemoryController.scala 100:37]
  reg  myID; // @[WriteMemoryController.scala 106:21]
  reg [31:0] _RAND_9;
  reg  isWrite; // @[WriteMemoryController.scala 108:24]
  reg [31:0] _RAND_10;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire [19:0] _T_10; // @[WriteMemoryController.scala 121:44]
  wire [21:0] _T_11; // @[WriteMemoryController.scala 121:69]
  wire  _T_12; // @[helpers.scala 27:24]
  wire  _T_13; // @[helpers.scala 27:47]
  wire  _T_14; // @[helpers.scala 27:40]
  wire  _T_16; // @[helpers.scala 28:15]
  wire  _T_17; // @[helpers.scala 28:38]
  wire  _T_18; // @[helpers.scala 28:31]
  wire  _T_20; // @[helpers.scala 29:17]
  wire  _T_21; // @[helpers.scala 29:40]
  wire  _T_22; // @[helpers.scala 29:33]
  wire [1:0] _T_28; // @[helpers.scala 39:32]
  wire [4:0] _T_29; // @[Cat.scala 29:58]
  wire [7:0] _T_43; // @[helpers.scala 50:12]
  wire [7:0] _T_44; // @[helpers.scala 49:10]
  wire [7:0] _T_45; // @[helpers.scala 48:19]
  wire [10:0] _GEN_31; // @[helpers.scala 20:26]
  wire [10:0] _T_47; // @[helpers.scala 20:26]
  wire [62:0] _GEN_32; // @[WriteMemoryController.scala 127:41]
  wire [62:0] _T_50; // @[WriteMemoryController.scala 127:41]
  wire [63:0] _T_52;
  wire [31:0] _T_53; // @[WriteMemoryController.scala 127:121]
  wire [31:0] _T_54; // @[WriteMemoryController.scala 127:121]
  wire [10:0] _GEN_10; // @[WriteMemoryController.scala 117:28]
  wire  _T_55; // @[WriteMemoryController.scala 139:15]
  wire  _T_56; // @[WriteMemoryController.scala 139:47]
  wire  _T_57; // @[WriteMemoryController.scala 139:30]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire [3:0] _T_59; // @[WriteMemoryController.scala 144:36]
  wire  _T_61; // @[WriteMemoryController.scala 146:18]
  wire [10:0] _GEN_14; // @[WriteMemoryController.scala 142:29]
  wire [10:0] _GEN_18; // @[WriteMemoryController.scala 139:76]
  wire  _T_62; // @[WriteMemoryController.scala 156:15]
  wire  _T_64; // @[WriteMemoryController.scala 156:32]
  wire  _T_65; // @[WriteMemoryController.scala 158:27]
  wire  _T_68; // @[Decoupled.scala 40:37]
  assign _T_4 = state == 2'h3; // @[WriteMemoryController.scala 89:21]
  assign _T_5 = {ptr,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_29 = {{29'd0}, _T_5}; // @[WriteMemoryController.scala 100:37]
  assign _T_9 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_NodeReq_bits_address[21:2]; // @[WriteMemoryController.scala 121:44]
  assign _T_11 = {_T_10, 2'h0}; // @[WriteMemoryController.scala 121:69]
  assign _T_12 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_13 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_14 = _T_12 | _T_13; // @[helpers.scala 27:40]
  assign _T_16 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_17 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_18 = _T_16 | _T_17; // @[helpers.scala 28:31]
  assign _T_20 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_21 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_22 = _T_20 | _T_21; // @[helpers.scala 29:33]
  assign _T_28 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_29 = {_T_28,3'h0}; // @[Cat.scala 29:58]
  assign _T_43 = _T_22 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_44 = _T_18 ? 8'h1 : _T_43; // @[helpers.scala 49:10]
  assign _T_45 = _T_14 ? 8'h3 : _T_44; // @[helpers.scala 48:19]
  assign _GEN_31 = {{3'd0}, _T_45}; // @[helpers.scala 20:26]
  assign _T_47 = _GEN_31 << _T_28; // @[helpers.scala 20:26]
  assign _GEN_32 = {{31'd0}, io_NodeReq_bits_data}; // @[WriteMemoryController.scala 127:41]
  assign _T_50 = _GEN_32 << _T_29; // @[WriteMemoryController.scala 127:41]
  assign _T_52 = {{1'd0}, _T_50};
  assign _T_53 = _T_52[31:0]; // @[WriteMemoryController.scala 127:121]
  assign _T_54 = _T_52[63:32]; // @[WriteMemoryController.scala 127:121]
  assign _GEN_10 = _T_9 ? _T_47 : {{3'd0}, sendbytemask}; // @[WriteMemoryController.scala 117:28]
  assign _T_55 = state == 2'h1; // @[WriteMemoryController.scala 139:15]
  assign _T_56 = sendbytemask != 8'h0; // @[WriteMemoryController.scala 139:47]
  assign _T_57 = _T_55 & _T_56; // @[WriteMemoryController.scala 139:30]
  assign _T_58 = io_MemReq_ready & io_MemReq_valid; // @[Decoupled.scala 40:37]
  assign _T_59 = sendbytemask[7:4]; // @[WriteMemoryController.scala 144:36]
  assign _T_61 = ptr + 1'h1; // @[WriteMemoryController.scala 146:18]
  assign _GEN_14 = _T_58 ? {{7'd0}, _T_59} : _GEN_10; // @[WriteMemoryController.scala 142:29]
  assign _GEN_18 = _T_57 ? _GEN_14 : _GEN_10; // @[WriteMemoryController.scala 139:76]
  assign _T_62 = state == 2'h2; // @[WriteMemoryController.scala 156:15]
  assign _T_64 = _T_62 & io_MemResp_valid; // @[WriteMemoryController.scala 156:32]
  assign _T_65 = sendbytemask == 8'h0; // @[WriteMemoryController.scala 158:27]
  assign _T_68 = io_output_ready & io_output_valid; // @[Decoupled.scala 40:37]
  assign io_NodeReq_ready = state == 2'h0; // @[WriteMemoryController.scala 87:20]
  assign io_MemReq_valid = _T_55 & _T_56; // @[WriteMemoryController.scala 99:19 WriteMemoryController.scala 140:21]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_29; // @[WriteMemoryController.scala 100:23]
  assign io_MemReq_bits_data = ptr ? linebuffer_1 : linebuffer_0; // @[WriteMemoryController.scala 102:23]
  assign io_MemReq_bits_mask = sendbytemask[3:0]; // @[WriteMemoryController.scala 103:23]
  assign io_MemReq_bits_tag = {{7'd0}, myID}; // @[WriteMemoryController.scala 107:22]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[WriteMemoryController.scala 110:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[WriteMemoryController.scala 109:26]
  assign io_output_valid = state == 2'h3; // @[WriteMemoryController.scala 95:19 WriteMemoryController.scala 168:21]
  assign io_output_bits_RouteID = request_R_RouteID; // @[WriteMemoryController.scala 98:26]
  assign io_free = state == 2'h0; // @[WriteMemoryController.scala 85:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ID = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_RouteID = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  request_R_taskID = _RAND_2[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  sendbytemask = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ReqAddress = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ptr = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  linebuffer_0 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  linebuffer_1 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  myID = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  isWrite = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    ID <= reset | ID;
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_9) begin
        request_R_RouteID <= io_NodeReq_bits_RouteID;
      end
    end
    if (reset) begin
      request_R_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_18[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_9) begin
        ReqAddress <= {{10'd0}, _T_11};
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (_T_4) begin
        ptr <= 1'h0;
      end else begin
        if (_T_57) begin
          if (_T_58) begin
            ptr <= _T_61;
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (_T_9) begin
        linebuffer_0 <= _T_53;
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (_T_9) begin
        linebuffer_1 <= _T_54;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_4) begin
        if (_T_68) begin
          state <= 2'h0;
        end else begin
          if (_T_64) begin
            if (_T_65) begin
              state <= 2'h3;
            end else begin
              state <= 2'h1;
            end
          end else begin
            if (_T_57) begin
              if (_T_58) begin
                state <= 2'h2;
              end else begin
                if (_T_9) begin
                  state <= 2'h1;
                end
              end
            end else begin
              if (_T_9) begin
                state <= 2'h1;
              end
            end
          end
        end
      end else begin
        if (_T_64) begin
          if (_T_65) begin
            state <= 2'h3;
          end else begin
            state <= 2'h1;
          end
        end else begin
          if (_T_57) begin
            if (_T_58) begin
              state <= 2'h2;
            end else begin
              if (_T_9) begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_9) begin
              state <= 2'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      myID <= 1'h0;
    end else begin
      myID <= ID;
    end
    if (reset) begin
      isWrite <= 1'h0;
    end else begin
      isWrite <= 1'h1;
    end
  end
endmodule
module WriteMemoryController(
  input         clock,
  input         reset,
  output        io_WriteIn_0_ready,
  input         io_WriteIn_0_valid,
  input  [21:0] io_WriteIn_0_bits_address,
  input  [31:0] io_WriteIn_0_bits_data,
  input  [4:0]  io_WriteIn_0_bits_taskID,
  output        io_WriteIn_1_ready,
  input         io_WriteIn_1_valid,
  input  [21:0] io_WriteIn_1_bits_address,
  input  [31:0] io_WriteIn_1_bits_data,
  input  [4:0]  io_WriteIn_1_bits_taskID,
  output        io_WriteIn_2_ready,
  input         io_WriteIn_2_valid,
  input  [21:0] io_WriteIn_2_bits_address,
  input  [31:0] io_WriteIn_2_bits_data,
  input  [4:0]  io_WriteIn_2_bits_taskID,
  output        io_WriteIn_3_ready,
  input         io_WriteIn_3_valid,
  input  [21:0] io_WriteIn_3_bits_address,
  input  [31:0] io_WriteIn_3_bits_data,
  input  [4:0]  io_WriteIn_3_bits_taskID,
  output        io_WriteIn_4_ready,
  input         io_WriteIn_4_valid,
  input  [21:0] io_WriteIn_4_bits_address,
  input  [31:0] io_WriteIn_4_bits_data,
  input  [4:0]  io_WriteIn_4_bits_taskID,
  output        io_WriteIn_5_ready,
  input         io_WriteIn_5_valid,
  input  [21:0] io_WriteIn_5_bits_address,
  input  [31:0] io_WriteIn_5_bits_data,
  input  [4:0]  io_WriteIn_5_bits_taskID,
  output        io_WriteIn_6_ready,
  input         io_WriteIn_6_valid,
  input  [21:0] io_WriteIn_6_bits_address,
  input  [31:0] io_WriteIn_6_bits_data,
  input  [4:0]  io_WriteIn_6_bits_taskID,
  output        io_WriteIn_7_ready,
  input         io_WriteIn_7_valid,
  input  [21:0] io_WriteIn_7_bits_address,
  input  [31:0] io_WriteIn_7_bits_data,
  input  [4:0]  io_WriteIn_7_bits_taskID,
  output        io_WriteIn_8_ready,
  input         io_WriteIn_8_valid,
  input  [21:0] io_WriteIn_8_bits_address,
  input  [31:0] io_WriteIn_8_bits_data,
  input  [4:0]  io_WriteIn_8_bits_taskID,
  output        io_WriteOut_0_valid,
  output        io_WriteOut_1_valid,
  output        io_WriteOut_2_valid,
  output        io_WriteOut_3_valid,
  output        io_WriteOut_4_valid,
  output        io_WriteOut_5_valid,
  output        io_WriteOut_6_valid,
  output        io_WriteOut_7_valid,
  output        io_WriteOut_8_valid,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag
);
  wire  in_arb_clock; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_0_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_0_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_0_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_0_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_0_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_1_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_1_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_1_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_1_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_1_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_2_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_2_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_2_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_2_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_2_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_3_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_3_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_3_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_3_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_3_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_4_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_4_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_4_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_4_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_4_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_5_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_5_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_5_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_5_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_5_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_6_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_6_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_6_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_6_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_6_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_7_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_7_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_7_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_7_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_7_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_8_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_in_8_valid; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_in_8_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_in_8_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_in_8_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_out_ready; // @[WriteMemoryController.scala 194:25]
  wire  in_arb_io_out_valid; // @[WriteMemoryController.scala 194:25]
  wire [15:0] in_arb_io_out_bits_RouteID; // @[WriteMemoryController.scala 194:25]
  wire [21:0] in_arb_io_out_bits_address; // @[WriteMemoryController.scala 194:25]
  wire [31:0] in_arb_io_out_bits_data; // @[WriteMemoryController.scala 194:25]
  wire [4:0] in_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 194:25]
  wire [7:0] in_arb_io_out_bits_Typ; // @[WriteMemoryController.scala 194:25]
  wire  alloc_arb_io_in_0_ready; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_in_0_valid; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_in_1_ready; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_in_1_valid; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_out_ready; // @[WriteMemoryController.scala 196:25]
  wire  alloc_arb_io_out_valid; // @[WriteMemoryController.scala 196:25]
  wire  cachereq_arb_io_in_0_ready; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_0_valid; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_0_bits_addr; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_0_bits_data; // @[WriteMemoryController.scala 199:31]
  wire [3:0] cachereq_arb_io_in_0_bits_mask; // @[WriteMemoryController.scala 199:31]
  wire [7:0] cachereq_arb_io_in_0_bits_tag; // @[WriteMemoryController.scala 199:31]
  wire [4:0] cachereq_arb_io_in_0_bits_taskID; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_0_bits_iswrite; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_1_ready; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_1_valid; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_1_bits_addr; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_in_1_bits_data; // @[WriteMemoryController.scala 199:31]
  wire [3:0] cachereq_arb_io_in_1_bits_mask; // @[WriteMemoryController.scala 199:31]
  wire [7:0] cachereq_arb_io_in_1_bits_tag; // @[WriteMemoryController.scala 199:31]
  wire [4:0] cachereq_arb_io_in_1_bits_taskID; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_in_1_bits_iswrite; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_out_ready; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_out_valid; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_out_bits_addr; // @[WriteMemoryController.scala 199:31]
  wire [31:0] cachereq_arb_io_out_bits_data; // @[WriteMemoryController.scala 199:31]
  wire [3:0] cachereq_arb_io_out_bits_mask; // @[WriteMemoryController.scala 199:31]
  wire [7:0] cachereq_arb_io_out_bits_tag; // @[WriteMemoryController.scala 199:31]
  wire [4:0] cachereq_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 199:31]
  wire  cachereq_arb_io_out_bits_iswrite; // @[WriteMemoryController.scala 199:31]
  wire  cacheresp_demux_io_en; // @[WriteMemoryController.scala 201:31]
  wire [31:0] cacheresp_demux_io_input_data; // @[WriteMemoryController.scala 201:31]
  wire [7:0] cacheresp_demux_io_input_tag; // @[WriteMemoryController.scala 201:31]
  wire  cacheresp_demux_io_sel; // @[WriteMemoryController.scala 201:31]
  wire  cacheresp_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 201:31]
  wire [31:0] cacheresp_demux_io_outputs_0_data; // @[WriteMemoryController.scala 201:31]
  wire [7:0] cacheresp_demux_io_outputs_0_tag; // @[WriteMemoryController.scala 201:31]
  wire  cacheresp_demux_io_outputs_1_valid; // @[WriteMemoryController.scala 201:31]
  wire [31:0] cacheresp_demux_io_outputs_1_data; // @[WriteMemoryController.scala 201:31]
  wire [7:0] cacheresp_demux_io_outputs_1_tag; // @[WriteMemoryController.scala 201:31]
  wire  out_arb_clock; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_0_ready; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_0_valid; // @[WriteMemoryController.scala 204:25]
  wire [15:0] out_arb_io_in_0_bits_RouteID; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_1_ready; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_in_1_valid; // @[WriteMemoryController.scala 204:25]
  wire [15:0] out_arb_io_in_1_bits_RouteID; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_out_ready; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_out_valid; // @[WriteMemoryController.scala 204:25]
  wire [15:0] out_arb_io_out_bits_RouteID; // @[WriteMemoryController.scala 204:25]
  wire  out_arb_io_chosen; // @[WriteMemoryController.scala 204:25]
  wire  out_demux_clock; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_reset; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_outputs_1_valid; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_outputs_2_valid; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_outputs_3_valid; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_outputs_4_valid; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_outputs_5_valid; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_outputs_6_valid; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_outputs_7_valid; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_outputs_8_valid; // @[WriteMemoryController.scala 205:25]
  wire [15:0] out_demux_io_input_RouteID; // @[WriteMemoryController.scala 205:25]
  wire  out_demux_io_enable; // @[WriteMemoryController.scala 205:25]
  wire  WriteTable_0_clock; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_reset; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_NodeReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_NodeReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [15:0] WriteTable_0_io_NodeReq_bits_RouteID; // @[WriteMemoryController.scala 223:29]
  wire [21:0] WriteTable_0_io_NodeReq_bits_address; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_0_io_NodeReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [4:0] WriteTable_0_io_NodeReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire [7:0] WriteTable_0_io_NodeReq_bits_Typ; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_0_io_MemReq_bits_addr; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_0_io_MemReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [3:0] WriteTable_0_io_MemReq_bits_mask; // @[WriteMemoryController.scala 223:29]
  wire [4:0] WriteTable_0_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_MemResp_valid; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_output_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_output_valid; // @[WriteMemoryController.scala 223:29]
  wire [15:0] WriteTable_0_io_output_bits_RouteID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_0_io_free; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_clock; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_reset; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_NodeReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_NodeReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [15:0] WriteTable_1_io_NodeReq_bits_RouteID; // @[WriteMemoryController.scala 223:29]
  wire [21:0] WriteTable_1_io_NodeReq_bits_address; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_1_io_NodeReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [4:0] WriteTable_1_io_NodeReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire [7:0] WriteTable_1_io_NodeReq_bits_Typ; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemReq_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemReq_valid; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_1_io_MemReq_bits_addr; // @[WriteMemoryController.scala 223:29]
  wire [31:0] WriteTable_1_io_MemReq_bits_data; // @[WriteMemoryController.scala 223:29]
  wire [3:0] WriteTable_1_io_MemReq_bits_mask; // @[WriteMemoryController.scala 223:29]
  wire [7:0] WriteTable_1_io_MemReq_bits_tag; // @[WriteMemoryController.scala 223:29]
  wire [4:0] WriteTable_1_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_MemResp_valid; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_output_ready; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_output_valid; // @[WriteMemoryController.scala 223:29]
  wire [15:0] WriteTable_1_io_output_bits_RouteID; // @[WriteMemoryController.scala 223:29]
  wire  WriteTable_1_io_free; // @[WriteMemoryController.scala 223:29]
  ArbiterTree in_arb ( // @[WriteMemoryController.scala 194:25]
    .clock(in_arb_clock),
    .io_in_0_ready(in_arb_io_in_0_ready),
    .io_in_0_valid(in_arb_io_in_0_valid),
    .io_in_0_bits_address(in_arb_io_in_0_bits_address),
    .io_in_0_bits_data(in_arb_io_in_0_bits_data),
    .io_in_0_bits_taskID(in_arb_io_in_0_bits_taskID),
    .io_in_1_ready(in_arb_io_in_1_ready),
    .io_in_1_valid(in_arb_io_in_1_valid),
    .io_in_1_bits_address(in_arb_io_in_1_bits_address),
    .io_in_1_bits_data(in_arb_io_in_1_bits_data),
    .io_in_1_bits_taskID(in_arb_io_in_1_bits_taskID),
    .io_in_2_ready(in_arb_io_in_2_ready),
    .io_in_2_valid(in_arb_io_in_2_valid),
    .io_in_2_bits_address(in_arb_io_in_2_bits_address),
    .io_in_2_bits_data(in_arb_io_in_2_bits_data),
    .io_in_2_bits_taskID(in_arb_io_in_2_bits_taskID),
    .io_in_3_ready(in_arb_io_in_3_ready),
    .io_in_3_valid(in_arb_io_in_3_valid),
    .io_in_3_bits_address(in_arb_io_in_3_bits_address),
    .io_in_3_bits_data(in_arb_io_in_3_bits_data),
    .io_in_3_bits_taskID(in_arb_io_in_3_bits_taskID),
    .io_in_4_ready(in_arb_io_in_4_ready),
    .io_in_4_valid(in_arb_io_in_4_valid),
    .io_in_4_bits_address(in_arb_io_in_4_bits_address),
    .io_in_4_bits_data(in_arb_io_in_4_bits_data),
    .io_in_4_bits_taskID(in_arb_io_in_4_bits_taskID),
    .io_in_5_ready(in_arb_io_in_5_ready),
    .io_in_5_valid(in_arb_io_in_5_valid),
    .io_in_5_bits_address(in_arb_io_in_5_bits_address),
    .io_in_5_bits_data(in_arb_io_in_5_bits_data),
    .io_in_5_bits_taskID(in_arb_io_in_5_bits_taskID),
    .io_in_6_ready(in_arb_io_in_6_ready),
    .io_in_6_valid(in_arb_io_in_6_valid),
    .io_in_6_bits_address(in_arb_io_in_6_bits_address),
    .io_in_6_bits_data(in_arb_io_in_6_bits_data),
    .io_in_6_bits_taskID(in_arb_io_in_6_bits_taskID),
    .io_in_7_ready(in_arb_io_in_7_ready),
    .io_in_7_valid(in_arb_io_in_7_valid),
    .io_in_7_bits_address(in_arb_io_in_7_bits_address),
    .io_in_7_bits_data(in_arb_io_in_7_bits_data),
    .io_in_7_bits_taskID(in_arb_io_in_7_bits_taskID),
    .io_in_8_ready(in_arb_io_in_8_ready),
    .io_in_8_valid(in_arb_io_in_8_valid),
    .io_in_8_bits_address(in_arb_io_in_8_bits_address),
    .io_in_8_bits_data(in_arb_io_in_8_bits_data),
    .io_in_8_bits_taskID(in_arb_io_in_8_bits_taskID),
    .io_out_ready(in_arb_io_out_ready),
    .io_out_valid(in_arb_io_out_valid),
    .io_out_bits_RouteID(in_arb_io_out_bits_RouteID),
    .io_out_bits_address(in_arb_io_out_bits_address),
    .io_out_bits_data(in_arb_io_out_bits_data),
    .io_out_bits_taskID(in_arb_io_out_bits_taskID),
    .io_out_bits_Typ(in_arb_io_out_bits_Typ)
  );
  Arbiter alloc_arb ( // @[WriteMemoryController.scala 196:25]
    .io_in_0_ready(alloc_arb_io_in_0_ready),
    .io_in_0_valid(alloc_arb_io_in_0_valid),
    .io_in_1_ready(alloc_arb_io_in_1_ready),
    .io_in_1_valid(alloc_arb_io_in_1_valid),
    .io_out_ready(alloc_arb_io_out_ready),
    .io_out_valid(alloc_arb_io_out_valid)
  );
  Arbiter_1 cachereq_arb ( // @[WriteMemoryController.scala 199:31]
    .io_in_0_ready(cachereq_arb_io_in_0_ready),
    .io_in_0_valid(cachereq_arb_io_in_0_valid),
    .io_in_0_bits_addr(cachereq_arb_io_in_0_bits_addr),
    .io_in_0_bits_data(cachereq_arb_io_in_0_bits_data),
    .io_in_0_bits_mask(cachereq_arb_io_in_0_bits_mask),
    .io_in_0_bits_tag(cachereq_arb_io_in_0_bits_tag),
    .io_in_0_bits_taskID(cachereq_arb_io_in_0_bits_taskID),
    .io_in_0_bits_iswrite(cachereq_arb_io_in_0_bits_iswrite),
    .io_in_1_ready(cachereq_arb_io_in_1_ready),
    .io_in_1_valid(cachereq_arb_io_in_1_valid),
    .io_in_1_bits_addr(cachereq_arb_io_in_1_bits_addr),
    .io_in_1_bits_data(cachereq_arb_io_in_1_bits_data),
    .io_in_1_bits_mask(cachereq_arb_io_in_1_bits_mask),
    .io_in_1_bits_tag(cachereq_arb_io_in_1_bits_tag),
    .io_in_1_bits_taskID(cachereq_arb_io_in_1_bits_taskID),
    .io_in_1_bits_iswrite(cachereq_arb_io_in_1_bits_iswrite),
    .io_out_ready(cachereq_arb_io_out_ready),
    .io_out_valid(cachereq_arb_io_out_valid),
    .io_out_bits_addr(cachereq_arb_io_out_bits_addr),
    .io_out_bits_data(cachereq_arb_io_out_bits_data),
    .io_out_bits_mask(cachereq_arb_io_out_bits_mask),
    .io_out_bits_tag(cachereq_arb_io_out_bits_tag),
    .io_out_bits_taskID(cachereq_arb_io_out_bits_taskID),
    .io_out_bits_iswrite(cachereq_arb_io_out_bits_iswrite)
  );
  Demux cacheresp_demux ( // @[WriteMemoryController.scala 201:31]
    .io_en(cacheresp_demux_io_en),
    .io_input_data(cacheresp_demux_io_input_data),
    .io_input_tag(cacheresp_demux_io_input_tag),
    .io_sel(cacheresp_demux_io_sel),
    .io_outputs_0_valid(cacheresp_demux_io_outputs_0_valid),
    .io_outputs_0_data(cacheresp_demux_io_outputs_0_data),
    .io_outputs_0_tag(cacheresp_demux_io_outputs_0_tag),
    .io_outputs_1_valid(cacheresp_demux_io_outputs_1_valid),
    .io_outputs_1_data(cacheresp_demux_io_outputs_1_data),
    .io_outputs_1_tag(cacheresp_demux_io_outputs_1_tag)
  );
  RRArbiter out_arb ( // @[WriteMemoryController.scala 204:25]
    .clock(out_arb_clock),
    .io_in_0_ready(out_arb_io_in_0_ready),
    .io_in_0_valid(out_arb_io_in_0_valid),
    .io_in_0_bits_RouteID(out_arb_io_in_0_bits_RouteID),
    .io_in_1_ready(out_arb_io_in_1_ready),
    .io_in_1_valid(out_arb_io_in_1_valid),
    .io_in_1_bits_RouteID(out_arb_io_in_1_bits_RouteID),
    .io_out_ready(out_arb_io_out_ready),
    .io_out_valid(out_arb_io_out_valid),
    .io_out_bits_RouteID(out_arb_io_out_bits_RouteID),
    .io_chosen(out_arb_io_chosen)
  );
  DeMuxTree out_demux ( // @[WriteMemoryController.scala 205:25]
    .clock(out_demux_clock),
    .reset(out_demux_reset),
    .io_outputs_0_valid(out_demux_io_outputs_0_valid),
    .io_outputs_1_valid(out_demux_io_outputs_1_valid),
    .io_outputs_2_valid(out_demux_io_outputs_2_valid),
    .io_outputs_3_valid(out_demux_io_outputs_3_valid),
    .io_outputs_4_valid(out_demux_io_outputs_4_valid),
    .io_outputs_5_valid(out_demux_io_outputs_5_valid),
    .io_outputs_6_valid(out_demux_io_outputs_6_valid),
    .io_outputs_7_valid(out_demux_io_outputs_7_valid),
    .io_outputs_8_valid(out_demux_io_outputs_8_valid),
    .io_input_RouteID(out_demux_io_input_RouteID),
    .io_enable(out_demux_io_enable)
  );
  WriteTableEntry WriteTable_0 ( // @[WriteMemoryController.scala 223:29]
    .clock(WriteTable_0_clock),
    .reset(WriteTable_0_reset),
    .io_NodeReq_ready(WriteTable_0_io_NodeReq_ready),
    .io_NodeReq_valid(WriteTable_0_io_NodeReq_valid),
    .io_NodeReq_bits_RouteID(WriteTable_0_io_NodeReq_bits_RouteID),
    .io_NodeReq_bits_address(WriteTable_0_io_NodeReq_bits_address),
    .io_NodeReq_bits_data(WriteTable_0_io_NodeReq_bits_data),
    .io_NodeReq_bits_taskID(WriteTable_0_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(WriteTable_0_io_NodeReq_bits_Typ),
    .io_MemReq_ready(WriteTable_0_io_MemReq_ready),
    .io_MemReq_valid(WriteTable_0_io_MemReq_valid),
    .io_MemReq_bits_addr(WriteTable_0_io_MemReq_bits_addr),
    .io_MemReq_bits_data(WriteTable_0_io_MemReq_bits_data),
    .io_MemReq_bits_mask(WriteTable_0_io_MemReq_bits_mask),
    .io_MemReq_bits_taskID(WriteTable_0_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(WriteTable_0_io_MemReq_bits_iswrite),
    .io_MemResp_valid(WriteTable_0_io_MemResp_valid),
    .io_output_ready(WriteTable_0_io_output_ready),
    .io_output_valid(WriteTable_0_io_output_valid),
    .io_output_bits_RouteID(WriteTable_0_io_output_bits_RouteID),
    .io_free(WriteTable_0_io_free)
  );
  WriteTableEntry_1 WriteTable_1 ( // @[WriteMemoryController.scala 223:29]
    .clock(WriteTable_1_clock),
    .reset(WriteTable_1_reset),
    .io_NodeReq_ready(WriteTable_1_io_NodeReq_ready),
    .io_NodeReq_valid(WriteTable_1_io_NodeReq_valid),
    .io_NodeReq_bits_RouteID(WriteTable_1_io_NodeReq_bits_RouteID),
    .io_NodeReq_bits_address(WriteTable_1_io_NodeReq_bits_address),
    .io_NodeReq_bits_data(WriteTable_1_io_NodeReq_bits_data),
    .io_NodeReq_bits_taskID(WriteTable_1_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(WriteTable_1_io_NodeReq_bits_Typ),
    .io_MemReq_ready(WriteTable_1_io_MemReq_ready),
    .io_MemReq_valid(WriteTable_1_io_MemReq_valid),
    .io_MemReq_bits_addr(WriteTable_1_io_MemReq_bits_addr),
    .io_MemReq_bits_data(WriteTable_1_io_MemReq_bits_data),
    .io_MemReq_bits_mask(WriteTable_1_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(WriteTable_1_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(WriteTable_1_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(WriteTable_1_io_MemReq_bits_iswrite),
    .io_MemResp_valid(WriteTable_1_io_MemResp_valid),
    .io_output_ready(WriteTable_1_io_output_ready),
    .io_output_valid(WriteTable_1_io_output_valid),
    .io_output_bits_RouteID(WriteTable_1_io_output_bits_RouteID),
    .io_free(WriteTable_1_io_free)
  );
  assign io_WriteIn_0_ready = in_arb_io_in_0_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteIn_1_ready = in_arb_io_in_1_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteIn_2_ready = in_arb_io_in_2_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteIn_3_ready = in_arb_io_in_3_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteIn_4_ready = in_arb_io_in_4_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteIn_5_ready = in_arb_io_in_5_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteIn_6_ready = in_arb_io_in_6_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteIn_7_ready = in_arb_io_in_7_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteIn_8_ready = in_arb_io_in_8_ready; // @[WriteMemoryController.scala 213:21]
  assign io_WriteOut_0_valid = out_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 214:20]
  assign io_WriteOut_1_valid = out_demux_io_outputs_1_valid; // @[WriteMemoryController.scala 214:20]
  assign io_WriteOut_2_valid = out_demux_io_outputs_2_valid; // @[WriteMemoryController.scala 214:20]
  assign io_WriteOut_3_valid = out_demux_io_outputs_3_valid; // @[WriteMemoryController.scala 214:20]
  assign io_WriteOut_4_valid = out_demux_io_outputs_4_valid; // @[WriteMemoryController.scala 214:20]
  assign io_WriteOut_5_valid = out_demux_io_outputs_5_valid; // @[WriteMemoryController.scala 214:20]
  assign io_WriteOut_6_valid = out_demux_io_outputs_6_valid; // @[WriteMemoryController.scala 214:20]
  assign io_WriteOut_7_valid = out_demux_io_outputs_7_valid; // @[WriteMemoryController.scala 214:20]
  assign io_WriteOut_8_valid = out_demux_io_outputs_8_valid; // @[WriteMemoryController.scala 214:20]
  assign io_MemReq_valid = cachereq_arb_io_out_valid; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_addr = cachereq_arb_io_out_bits_addr; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_data = cachereq_arb_io_out_bits_data; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_mask = cachereq_arb_io_out_bits_mask; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_tag = cachereq_arb_io_out_bits_tag; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_taskID = cachereq_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 261:13]
  assign io_MemReq_bits_iswrite = cachereq_arb_io_out_bits_iswrite; // @[WriteMemoryController.scala 261:13]
  assign in_arb_clock = clock;
  assign in_arb_io_in_0_valid = io_WriteIn_0_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_0_bits_address = io_WriteIn_0_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_0_bits_data = io_WriteIn_0_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_0_bits_taskID = io_WriteIn_0_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_1_valid = io_WriteIn_1_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_1_bits_address = io_WriteIn_1_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_1_bits_data = io_WriteIn_1_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_1_bits_taskID = io_WriteIn_1_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_2_valid = io_WriteIn_2_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_2_bits_address = io_WriteIn_2_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_2_bits_data = io_WriteIn_2_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_2_bits_taskID = io_WriteIn_2_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_3_valid = io_WriteIn_3_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_3_bits_address = io_WriteIn_3_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_3_bits_data = io_WriteIn_3_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_3_bits_taskID = io_WriteIn_3_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_4_valid = io_WriteIn_4_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_4_bits_address = io_WriteIn_4_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_4_bits_data = io_WriteIn_4_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_4_bits_taskID = io_WriteIn_4_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_5_valid = io_WriteIn_5_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_5_bits_address = io_WriteIn_5_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_5_bits_data = io_WriteIn_5_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_5_bits_taskID = io_WriteIn_5_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_6_valid = io_WriteIn_6_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_6_bits_address = io_WriteIn_6_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_6_bits_data = io_WriteIn_6_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_6_bits_taskID = io_WriteIn_6_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_7_valid = io_WriteIn_7_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_7_bits_address = io_WriteIn_7_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_7_bits_data = io_WriteIn_7_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_7_bits_taskID = io_WriteIn_7_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_8_valid = io_WriteIn_8_valid; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_8_bits_address = io_WriteIn_8_bits_address; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_8_bits_data = io_WriteIn_8_bits_data; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_in_8_bits_taskID = io_WriteIn_8_bits_taskID; // @[WriteMemoryController.scala 213:21]
  assign in_arb_io_out_ready = alloc_arb_io_out_valid; // @[WriteMemoryController.scala 256:23]
  assign alloc_arb_io_in_0_valid = WriteTable_0_io_free; // @[WriteMemoryController.scala 226:30]
  assign alloc_arb_io_in_1_valid = WriteTable_1_io_free; // @[WriteMemoryController.scala 226:30]
  assign alloc_arb_io_out_ready = in_arb_io_out_valid; // @[WriteMemoryController.scala 257:26]
  assign cachereq_arb_io_in_0_valid = WriteTable_0_io_MemReq_valid; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_addr = WriteTable_0_io_MemReq_bits_addr; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_data = WriteTable_0_io_MemReq_bits_data; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_mask = WriteTable_0_io_MemReq_bits_mask; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_tag = 8'h0; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_taskID = WriteTable_0_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_0_bits_iswrite = WriteTable_0_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_valid = WriteTable_1_io_MemReq_valid; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_addr = WriteTable_1_io_MemReq_bits_addr; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_data = WriteTable_1_io_MemReq_bits_data; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_mask = WriteTable_1_io_MemReq_bits_mask; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_tag = WriteTable_1_io_MemReq_bits_tag; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_taskID = WriteTable_1_io_MemReq_bits_taskID; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_in_1_bits_iswrite = WriteTable_1_io_MemReq_bits_iswrite; // @[WriteMemoryController.scala 232:27]
  assign cachereq_arb_io_out_ready = io_MemReq_ready; // @[WriteMemoryController.scala 261:13]
  assign cacheresp_demux_io_en = io_MemResp_valid; // @[WriteMemoryController.scala 264:25]
  assign cacheresp_demux_io_input_data = io_MemResp_bits_data; // @[WriteMemoryController.scala 265:28]
  assign cacheresp_demux_io_input_tag = io_MemResp_bits_tag; // @[WriteMemoryController.scala 265:28]
  assign cacheresp_demux_io_sel = io_MemResp_bits_tag[0]; // @[WriteMemoryController.scala 266:26]
  assign out_arb_clock = clock;
  assign out_arb_io_in_0_valid = WriteTable_0_io_output_valid; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_in_0_bits_RouteID = WriteTable_0_io_output_bits_RouteID; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_in_1_valid = WriteTable_1_io_output_valid; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_in_1_bits_RouteID = WriteTable_1_io_output_bits_RouteID; // @[WriteMemoryController.scala 238:22]
  assign out_arb_io_out_ready = 1'h1; // @[WriteMemoryController.scala 269:24]
  assign out_demux_clock = clock;
  assign out_demux_reset = reset;
  assign out_demux_io_input_RouteID = out_arb_io_out_bits_RouteID; // @[WriteMemoryController.scala 271:22]
  assign out_demux_io_enable = out_arb_io_out_ready & out_arb_io_out_valid; // @[WriteMemoryController.scala 270:23]
  assign WriteTable_0_clock = clock;
  assign WriteTable_0_reset = reset;
  assign WriteTable_0_io_NodeReq_valid = alloc_arb_io_in_0_ready & alloc_arb_io_in_0_valid; // @[WriteMemoryController.scala 228:34]
  assign WriteTable_0_io_NodeReq_bits_RouteID = in_arb_io_out_bits_RouteID; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_data = in_arb_io_out_bits_data; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_0_io_MemReq_ready = cachereq_arb_io_in_0_ready; // @[WriteMemoryController.scala 232:27]
  assign WriteTable_0_io_MemResp_valid = cacheresp_demux_io_outputs_0_valid; // @[WriteMemoryController.scala 235:28]
  assign WriteTable_0_io_output_ready = out_arb_io_in_0_ready; // @[WriteMemoryController.scala 238:22]
  assign WriteTable_1_clock = clock;
  assign WriteTable_1_reset = reset;
  assign WriteTable_1_io_NodeReq_valid = alloc_arb_io_in_1_ready & alloc_arb_io_in_1_valid; // @[WriteMemoryController.scala 228:34]
  assign WriteTable_1_io_NodeReq_bits_RouteID = in_arb_io_out_bits_RouteID; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_data = in_arb_io_out_bits_data; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[WriteMemoryController.scala 229:33]
  assign WriteTable_1_io_MemReq_ready = cachereq_arb_io_in_1_ready; // @[WriteMemoryController.scala 232:27]
  assign WriteTable_1_io_MemResp_valid = cacheresp_demux_io_outputs_1_valid; // @[WriteMemoryController.scala 235:28]
  assign WriteTable_1_io_output_ready = out_arb_io_in_1_ready; // @[WriteMemoryController.scala 238:22]
endmodule
module LockingRRArbiter_11(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [15:0] io_in_0_bits_RouteID,
  input  [31:0] io_in_0_bits_address,
  input  [4:0]  io_in_0_bits_taskID,
  input  [7:0]  io_in_0_bits_Typ,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [15:0] io_in_1_bits_RouteID,
  input  [31:0] io_in_1_bits_address,
  input  [4:0]  io_in_1_bits_taskID,
  input  [7:0]  io_in_1_bits_Typ,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [31:0] io_out_bits_address,
  output [4:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ,
  output        io_chosen
);
  wire  _T; // @[Decoupled.scala 40:37]
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Arbiter.scala 67:57]
  wire  _T_5; // @[Arbiter.scala 68:83]
  wire  _T_7; // @[Arbiter.scala 31:68]
  wire  _T_9; // @[Arbiter.scala 31:78]
  wire  _T_10; // @[Arbiter.scala 31:78]
  wire  _T_14; // @[Arbiter.scala 72:50]
  wire  _GEN_13; // @[Arbiter.scala 77:27]
  assign _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = 1'h1 > _T_1; // @[Arbiter.scala 67:57]
  assign _T_5 = io_in_1_valid & _T_3; // @[Arbiter.scala 68:83]
  assign _T_7 = _T_5 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_9 = _T_5 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_10 = _T_7 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_14 = _T_3 | _T_10; // @[Arbiter.scala 72:50]
  assign _GEN_13 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_9 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_14 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_RouteID = io_chosen ? io_in_1_bits_RouteID : io_in_0_bits_RouteID; // @[Arbiter.scala 42:15]
  assign io_out_bits_address = io_chosen ? io_in_1_bits_address : io_in_0_bits_address; // @[Arbiter.scala 42:15]
  assign io_out_bits_taskID = io_chosen ? io_in_1_bits_taskID : io_in_0_bits_taskID; // @[Arbiter.scala 42:15]
  assign io_out_bits_Typ = io_chosen ? io_in_1_bits_Typ : io_in_0_bits_Typ; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_5 | _GEN_13; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (_T) begin
      _T_1 <= io_chosen;
    end
  end
endmodule
module ArbiterTree_1(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_address,
  input  [4:0]  io_in_0_bits_taskID,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_address,
  input  [4:0]  io_in_1_bits_taskID,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_address,
  input  [4:0]  io_in_2_bits_taskID,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_address,
  input  [4:0]  io_in_3_bits_taskID,
  output        io_in_4_ready,
  input         io_in_4_valid,
  input  [31:0] io_in_4_bits_address,
  input  [4:0]  io_in_4_bits_taskID,
  output        io_in_5_ready,
  input         io_in_5_valid,
  input  [31:0] io_in_5_bits_address,
  input  [4:0]  io_in_5_bits_taskID,
  output        io_in_6_ready,
  input         io_in_6_valid,
  input  [31:0] io_in_6_bits_address,
  input  [4:0]  io_in_6_bits_taskID,
  output        io_in_7_ready,
  input         io_in_7_valid,
  input  [31:0] io_in_7_bits_address,
  input  [4:0]  io_in_7_bits_taskID,
  output        io_in_8_ready,
  input         io_in_8_valid,
  input  [31:0] io_in_8_bits_address,
  input  [4:0]  io_in_8_bits_taskID,
  output        io_in_9_ready,
  input         io_in_9_valid,
  input  [31:0] io_in_9_bits_address,
  input  [4:0]  io_in_9_bits_taskID,
  output        io_in_10_ready,
  input         io_in_10_valid,
  input  [31:0] io_in_10_bits_address,
  input  [4:0]  io_in_10_bits_taskID,
  output        io_in_11_ready,
  input         io_in_11_valid,
  input  [31:0] io_in_11_bits_address,
  input  [4:0]  io_in_11_bits_taskID,
  output        io_in_12_ready,
  input         io_in_12_valid,
  input  [31:0] io_in_12_bits_address,
  input  [4:0]  io_in_12_bits_taskID,
  output        io_in_13_ready,
  input         io_in_13_valid,
  input  [31:0] io_in_13_bits_address,
  input  [4:0]  io_in_13_bits_taskID,
  output        io_in_14_ready,
  input         io_in_14_valid,
  input  [31:0] io_in_14_bits_address,
  input  [4:0]  io_in_14_bits_taskID,
  output        io_in_15_ready,
  input         io_in_15_valid,
  input  [31:0] io_in_15_bits_address,
  input  [4:0]  io_in_15_bits_taskID,
  output        io_in_16_ready,
  input         io_in_16_valid,
  input  [31:0] io_in_16_bits_address,
  input  [4:0]  io_in_16_bits_taskID,
  output        io_in_17_ready,
  input         io_in_17_valid,
  input  [31:0] io_in_17_bits_address,
  input  [4:0]  io_in_17_bits_taskID,
  output        io_in_18_ready,
  input         io_in_18_valid,
  input  [31:0] io_in_18_bits_address,
  input  [4:0]  io_in_18_bits_taskID,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [31:0] io_out_bits_address,
  output [4:0]  io_out_bits_taskID,
  output [7:0]  io_out_bits_Typ
);
  wire  LockingRRArbiter_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_1_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_1_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_1_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_1_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_1_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_1_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_1_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_1_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_1_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_1_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_1_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_1_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_1_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_2_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_2_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_2_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_2_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_2_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_2_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_2_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_2_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_2_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_2_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_2_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_2_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_2_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_3_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_3_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_3_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_3_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_3_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_3_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_3_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_3_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_3_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_3_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_3_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_3_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_3_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_4_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_4_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_4_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_4_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_4_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_4_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_4_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_4_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_4_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_4_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_4_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_4_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_4_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_5_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_5_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_5_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_5_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_5_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_5_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_5_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_5_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_5_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_5_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_5_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_5_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_5_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_6_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_6_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_6_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_6_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_6_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_6_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_6_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_6_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_6_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_6_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_6_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_6_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_6_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_7_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_7_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_7_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_7_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_7_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_7_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_7_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_7_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_7_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_7_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_7_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_7_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_7_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_8_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_8_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_8_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_8_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_8_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_8_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_8_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_8_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_8_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_8_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_8_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_8_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_8_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_9_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_9_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_9_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_9_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_9_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_9_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_9_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_9_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_9_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_9_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_9_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_9_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_9_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_10_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_10_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_10_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_10_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_10_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_10_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_10_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_10_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_10_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_10_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_10_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_10_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_10_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_11_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_11_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_11_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_11_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_11_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_11_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_11_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_11_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_11_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_11_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_11_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_11_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_11_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_11_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_11_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_11_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_11_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_11_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_11_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_11_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_12_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_12_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_12_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_12_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_12_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_12_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_12_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_12_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_12_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_12_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_12_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_12_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_12_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_12_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_12_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_12_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_12_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_12_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_12_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_12_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_13_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_13_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_13_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_13_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_13_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_13_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_13_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_13_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_13_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_13_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_13_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_13_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_13_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_13_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_13_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_13_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_13_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_13_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_13_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_13_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_14_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_14_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_14_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_14_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_14_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_14_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_14_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_14_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_14_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_14_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_14_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_14_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_14_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_14_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_14_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_14_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_14_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_14_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_14_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_14_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_15_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_15_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_15_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_15_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_15_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_15_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_15_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_15_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_15_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_15_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_15_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_15_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_15_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_15_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_15_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_15_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_15_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_15_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_15_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_15_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_16_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_16_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_16_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_16_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_16_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_16_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_16_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_16_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_16_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_16_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_16_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_16_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_16_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_16_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_16_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_16_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_16_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_16_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_16_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_16_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_17_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_17_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_17_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_17_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_17_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_17_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_17_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_17_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_17_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_17_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_17_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_17_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_17_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_17_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_17_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_17_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_17_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_17_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_17_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_17_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_18_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_18_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_18_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_18_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_18_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_18_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_18_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_18_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_18_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_18_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_18_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_18_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_18_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_18_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_18_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_18_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_18_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_18_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_18_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_18_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_19_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_19_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_19_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_19_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_19_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_19_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_19_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_19_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_19_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_19_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_19_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_19_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_19_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_19_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_19_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_19_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_19_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_19_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_19_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_19_io_chosen; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_20_clock; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_20_io_in_0_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_20_io_in_0_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_20_io_in_0_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_20_io_in_0_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_20_io_in_0_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_20_io_in_0_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_20_io_in_1_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_20_io_in_1_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_20_io_in_1_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_20_io_in_1_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_20_io_in_1_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_20_io_in_1_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_20_io_out_ready; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_20_io_out_valid; // @[ArbiterTree.scala 32:13]
  wire [15:0] LockingRRArbiter_20_io_out_bits_RouteID; // @[ArbiterTree.scala 32:13]
  wire [31:0] LockingRRArbiter_20_io_out_bits_address; // @[ArbiterTree.scala 32:13]
  wire [4:0] LockingRRArbiter_20_io_out_bits_taskID; // @[ArbiterTree.scala 32:13]
  wire [7:0] LockingRRArbiter_20_io_out_bits_Typ; // @[ArbiterTree.scala 32:13]
  wire  LockingRRArbiter_20_io_chosen; // @[ArbiterTree.scala 32:13]
  LockingRRArbiter_11 LockingRRArbiter ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_clock),
    .io_in_0_ready(LockingRRArbiter_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_io_out_ready),
    .io_out_valid(LockingRRArbiter_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_1 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_1_clock),
    .io_in_0_ready(LockingRRArbiter_1_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_1_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_1_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_1_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_1_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_1_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_1_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_1_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_1_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_1_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_1_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_1_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_1_io_out_ready),
    .io_out_valid(LockingRRArbiter_1_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_1_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_1_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_1_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_1_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_1_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_2 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_2_clock),
    .io_in_0_ready(LockingRRArbiter_2_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_2_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_2_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_2_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_2_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_2_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_2_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_2_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_2_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_2_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_2_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_2_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_2_io_out_ready),
    .io_out_valid(LockingRRArbiter_2_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_2_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_2_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_2_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_2_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_2_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_3 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_3_clock),
    .io_in_0_ready(LockingRRArbiter_3_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_3_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_3_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_3_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_3_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_3_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_3_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_3_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_3_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_3_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_3_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_3_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_3_io_out_ready),
    .io_out_valid(LockingRRArbiter_3_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_3_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_3_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_3_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_3_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_3_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_4 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_4_clock),
    .io_in_0_ready(LockingRRArbiter_4_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_4_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_4_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_4_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_4_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_4_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_4_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_4_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_4_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_4_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_4_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_4_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_4_io_out_ready),
    .io_out_valid(LockingRRArbiter_4_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_4_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_4_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_4_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_4_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_4_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_5 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_5_clock),
    .io_in_0_ready(LockingRRArbiter_5_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_5_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_5_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_5_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_5_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_5_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_5_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_5_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_5_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_5_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_5_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_5_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_5_io_out_ready),
    .io_out_valid(LockingRRArbiter_5_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_5_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_5_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_5_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_5_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_5_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_6 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_6_clock),
    .io_in_0_ready(LockingRRArbiter_6_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_6_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_6_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_6_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_6_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_6_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_6_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_6_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_6_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_6_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_6_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_6_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_6_io_out_ready),
    .io_out_valid(LockingRRArbiter_6_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_6_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_6_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_6_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_6_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_6_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_7 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_7_clock),
    .io_in_0_ready(LockingRRArbiter_7_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_7_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_7_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_7_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_7_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_7_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_7_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_7_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_7_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_7_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_7_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_7_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_7_io_out_ready),
    .io_out_valid(LockingRRArbiter_7_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_7_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_7_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_7_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_7_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_7_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_8 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_8_clock),
    .io_in_0_ready(LockingRRArbiter_8_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_8_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_8_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_8_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_8_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_8_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_8_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_8_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_8_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_8_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_8_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_8_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_8_io_out_ready),
    .io_out_valid(LockingRRArbiter_8_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_8_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_8_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_8_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_8_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_8_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_9 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_9_clock),
    .io_in_0_ready(LockingRRArbiter_9_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_9_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_9_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_9_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_9_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_9_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_9_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_9_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_9_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_9_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_9_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_9_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_9_io_out_ready),
    .io_out_valid(LockingRRArbiter_9_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_9_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_9_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_9_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_9_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_9_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_10 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_10_clock),
    .io_in_0_ready(LockingRRArbiter_10_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_10_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_10_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_10_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_10_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_10_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_10_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_10_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_10_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_10_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_10_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_10_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_10_io_out_ready),
    .io_out_valid(LockingRRArbiter_10_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_10_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_10_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_10_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_10_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_10_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_11 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_11_clock),
    .io_in_0_ready(LockingRRArbiter_11_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_11_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_11_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_11_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_11_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_11_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_11_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_11_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_11_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_11_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_11_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_11_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_11_io_out_ready),
    .io_out_valid(LockingRRArbiter_11_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_11_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_11_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_11_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_11_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_11_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_12 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_12_clock),
    .io_in_0_ready(LockingRRArbiter_12_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_12_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_12_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_12_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_12_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_12_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_12_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_12_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_12_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_12_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_12_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_12_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_12_io_out_ready),
    .io_out_valid(LockingRRArbiter_12_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_12_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_12_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_12_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_12_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_12_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_13 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_13_clock),
    .io_in_0_ready(LockingRRArbiter_13_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_13_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_13_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_13_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_13_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_13_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_13_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_13_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_13_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_13_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_13_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_13_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_13_io_out_ready),
    .io_out_valid(LockingRRArbiter_13_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_13_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_13_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_13_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_13_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_13_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_14 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_14_clock),
    .io_in_0_ready(LockingRRArbiter_14_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_14_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_14_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_14_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_14_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_14_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_14_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_14_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_14_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_14_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_14_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_14_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_14_io_out_ready),
    .io_out_valid(LockingRRArbiter_14_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_14_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_14_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_14_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_14_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_14_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_15 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_15_clock),
    .io_in_0_ready(LockingRRArbiter_15_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_15_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_15_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_15_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_15_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_15_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_15_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_15_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_15_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_15_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_15_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_15_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_15_io_out_ready),
    .io_out_valid(LockingRRArbiter_15_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_15_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_15_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_15_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_15_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_15_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_16 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_16_clock),
    .io_in_0_ready(LockingRRArbiter_16_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_16_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_16_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_16_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_16_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_16_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_16_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_16_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_16_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_16_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_16_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_16_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_16_io_out_ready),
    .io_out_valid(LockingRRArbiter_16_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_16_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_16_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_16_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_16_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_16_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_17 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_17_clock),
    .io_in_0_ready(LockingRRArbiter_17_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_17_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_17_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_17_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_17_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_17_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_17_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_17_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_17_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_17_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_17_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_17_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_17_io_out_ready),
    .io_out_valid(LockingRRArbiter_17_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_17_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_17_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_17_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_17_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_17_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_18 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_18_clock),
    .io_in_0_ready(LockingRRArbiter_18_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_18_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_18_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_18_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_18_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_18_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_18_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_18_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_18_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_18_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_18_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_18_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_18_io_out_ready),
    .io_out_valid(LockingRRArbiter_18_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_18_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_18_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_18_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_18_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_18_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_19 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_19_clock),
    .io_in_0_ready(LockingRRArbiter_19_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_19_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_19_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_19_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_19_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_19_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_19_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_19_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_19_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_19_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_19_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_19_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_19_io_out_ready),
    .io_out_valid(LockingRRArbiter_19_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_19_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_19_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_19_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_19_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_19_io_chosen)
  );
  LockingRRArbiter_11 LockingRRArbiter_20 ( // @[ArbiterTree.scala 32:13]
    .clock(LockingRRArbiter_20_clock),
    .io_in_0_ready(LockingRRArbiter_20_io_in_0_ready),
    .io_in_0_valid(LockingRRArbiter_20_io_in_0_valid),
    .io_in_0_bits_RouteID(LockingRRArbiter_20_io_in_0_bits_RouteID),
    .io_in_0_bits_address(LockingRRArbiter_20_io_in_0_bits_address),
    .io_in_0_bits_taskID(LockingRRArbiter_20_io_in_0_bits_taskID),
    .io_in_0_bits_Typ(LockingRRArbiter_20_io_in_0_bits_Typ),
    .io_in_1_ready(LockingRRArbiter_20_io_in_1_ready),
    .io_in_1_valid(LockingRRArbiter_20_io_in_1_valid),
    .io_in_1_bits_RouteID(LockingRRArbiter_20_io_in_1_bits_RouteID),
    .io_in_1_bits_address(LockingRRArbiter_20_io_in_1_bits_address),
    .io_in_1_bits_taskID(LockingRRArbiter_20_io_in_1_bits_taskID),
    .io_in_1_bits_Typ(LockingRRArbiter_20_io_in_1_bits_Typ),
    .io_out_ready(LockingRRArbiter_20_io_out_ready),
    .io_out_valid(LockingRRArbiter_20_io_out_valid),
    .io_out_bits_RouteID(LockingRRArbiter_20_io_out_bits_RouteID),
    .io_out_bits_address(LockingRRArbiter_20_io_out_bits_address),
    .io_out_bits_taskID(LockingRRArbiter_20_io_out_bits_taskID),
    .io_out_bits_Typ(LockingRRArbiter_20_io_out_bits_Typ),
    .io_chosen(LockingRRArbiter_20_io_chosen)
  );
  assign io_in_0_ready = LockingRRArbiter_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_1_ready = LockingRRArbiter_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_2_ready = LockingRRArbiter_1_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_3_ready = LockingRRArbiter_1_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_4_ready = LockingRRArbiter_2_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_5_ready = LockingRRArbiter_2_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_6_ready = LockingRRArbiter_3_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_7_ready = LockingRRArbiter_3_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_8_ready = LockingRRArbiter_4_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_9_ready = LockingRRArbiter_4_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_10_ready = LockingRRArbiter_5_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_11_ready = LockingRRArbiter_5_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_12_ready = LockingRRArbiter_6_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_13_ready = LockingRRArbiter_6_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_14_ready = LockingRRArbiter_7_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_15_ready = LockingRRArbiter_7_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_16_ready = LockingRRArbiter_8_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_17_ready = LockingRRArbiter_8_io_in_1_ready; // @[ArbiterTree.scala 49:61]
  assign io_in_18_ready = LockingRRArbiter_9_io_in_0_ready; // @[ArbiterTree.scala 49:61]
  assign io_out_valid = LockingRRArbiter_20_io_out_valid; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_RouteID = LockingRRArbiter_20_io_out_bits_RouteID; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_address = LockingRRArbiter_20_io_out_bits_address; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_taskID = LockingRRArbiter_20_io_out_bits_taskID; // @[ArbiterTree.scala 65:12]
  assign io_out_bits_Typ = LockingRRArbiter_20_io_out_bits_Typ; // @[ArbiterTree.scala 65:12]
  assign LockingRRArbiter_clock = clock;
  assign LockingRRArbiter_io_in_0_valid = io_in_0_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_RouteID = 16'h0; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_address = io_in_0_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_taskID = io_in_0_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_valid = io_in_1_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_RouteID = 16'h1; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_address = io_in_1_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_taskID = io_in_1_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_io_out_ready = LockingRRArbiter_10_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_1_clock = clock;
  assign LockingRRArbiter_1_io_in_0_valid = io_in_2_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_RouteID = 16'h2; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_address = io_in_2_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_taskID = io_in_2_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_valid = io_in_3_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_bits_RouteID = 16'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_bits_address = io_in_3_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_bits_taskID = io_in_3_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_1_io_out_ready = LockingRRArbiter_10_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_2_clock = clock;
  assign LockingRRArbiter_2_io_in_0_valid = io_in_4_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_0_bits_RouteID = 16'h4; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_0_bits_address = io_in_4_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_0_bits_taskID = io_in_4_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_valid = io_in_5_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_bits_RouteID = 16'h5; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_bits_address = io_in_5_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_bits_taskID = io_in_5_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_2_io_out_ready = LockingRRArbiter_11_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_3_clock = clock;
  assign LockingRRArbiter_3_io_in_0_valid = io_in_6_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_0_bits_RouteID = 16'h6; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_0_bits_address = io_in_6_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_0_bits_taskID = io_in_6_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_valid = io_in_7_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_bits_RouteID = 16'h7; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_bits_address = io_in_7_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_bits_taskID = io_in_7_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_3_io_out_ready = LockingRRArbiter_11_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_4_clock = clock;
  assign LockingRRArbiter_4_io_in_0_valid = io_in_8_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_0_bits_RouteID = 16'h8; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_0_bits_address = io_in_8_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_0_bits_taskID = io_in_8_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_1_valid = io_in_9_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_1_bits_RouteID = 16'h9; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_1_bits_address = io_in_9_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_1_bits_taskID = io_in_9_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_4_io_out_ready = LockingRRArbiter_12_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_5_clock = clock;
  assign LockingRRArbiter_5_io_in_0_valid = io_in_10_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_in_0_bits_RouteID = 16'ha; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_in_0_bits_address = io_in_10_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_in_0_bits_taskID = io_in_10_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_in_1_valid = io_in_11_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_in_1_bits_RouteID = 16'hb; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_in_1_bits_address = io_in_11_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_in_1_bits_taskID = io_in_11_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_5_io_out_ready = LockingRRArbiter_12_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_6_clock = clock;
  assign LockingRRArbiter_6_io_in_0_valid = io_in_12_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_in_0_bits_RouteID = 16'hc; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_in_0_bits_address = io_in_12_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_in_0_bits_taskID = io_in_12_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_in_1_valid = io_in_13_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_in_1_bits_RouteID = 16'hd; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_in_1_bits_address = io_in_13_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_in_1_bits_taskID = io_in_13_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_6_io_out_ready = LockingRRArbiter_13_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_7_clock = clock;
  assign LockingRRArbiter_7_io_in_0_valid = io_in_14_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_in_0_bits_RouteID = 16'he; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_in_0_bits_address = io_in_14_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_in_0_bits_taskID = io_in_14_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_in_1_valid = io_in_15_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_in_1_bits_RouteID = 16'hf; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_in_1_bits_address = io_in_15_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_in_1_bits_taskID = io_in_15_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_7_io_out_ready = LockingRRArbiter_13_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_8_clock = clock;
  assign LockingRRArbiter_8_io_in_0_valid = io_in_16_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_in_0_bits_RouteID = 16'h10; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_in_0_bits_address = io_in_16_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_in_0_bits_taskID = io_in_16_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_in_1_valid = io_in_17_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_in_1_bits_RouteID = 16'h11; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_in_1_bits_address = io_in_17_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_in_1_bits_taskID = io_in_17_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_in_1_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_8_io_out_ready = LockingRRArbiter_14_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_9_clock = clock;
  assign LockingRRArbiter_9_io_in_0_valid = io_in_18_valid; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_9_io_in_0_bits_RouteID = 16'h12; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_9_io_in_0_bits_address = io_in_18_bits_address; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_9_io_in_0_bits_taskID = io_in_18_bits_taskID; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_9_io_in_0_bits_Typ = 8'h3; // @[ArbiterTree.scala 49:61]
  assign LockingRRArbiter_9_io_in_1_valid = 1'h0; // @[ArbiterTree.scala 52:67]
  assign LockingRRArbiter_9_io_in_1_bits_RouteID = 16'h0;
  assign LockingRRArbiter_9_io_in_1_bits_address = 32'h0;
  assign LockingRRArbiter_9_io_in_1_bits_taskID = 5'h0;
  assign LockingRRArbiter_9_io_in_1_bits_Typ = 8'h0;
  assign LockingRRArbiter_9_io_out_ready = LockingRRArbiter_14_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_clock = clock;
  assign LockingRRArbiter_10_io_in_0_valid = LockingRRArbiter_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_0_bits_RouteID = LockingRRArbiter_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_0_bits_address = LockingRRArbiter_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_0_bits_taskID = LockingRRArbiter_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_0_bits_Typ = LockingRRArbiter_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_valid = LockingRRArbiter_1_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_bits_RouteID = LockingRRArbiter_1_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_bits_address = LockingRRArbiter_1_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_bits_taskID = LockingRRArbiter_1_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_in_1_bits_Typ = LockingRRArbiter_1_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_10_io_out_ready = LockingRRArbiter_15_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_clock = clock;
  assign LockingRRArbiter_11_io_in_0_valid = LockingRRArbiter_2_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_in_0_bits_RouteID = LockingRRArbiter_2_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_in_0_bits_address = LockingRRArbiter_2_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_in_0_bits_taskID = LockingRRArbiter_2_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_in_0_bits_Typ = LockingRRArbiter_2_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_in_1_valid = LockingRRArbiter_3_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_in_1_bits_RouteID = LockingRRArbiter_3_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_in_1_bits_address = LockingRRArbiter_3_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_in_1_bits_taskID = LockingRRArbiter_3_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_in_1_bits_Typ = LockingRRArbiter_3_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_11_io_out_ready = LockingRRArbiter_15_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_clock = clock;
  assign LockingRRArbiter_12_io_in_0_valid = LockingRRArbiter_4_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_in_0_bits_RouteID = LockingRRArbiter_4_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_in_0_bits_address = LockingRRArbiter_4_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_in_0_bits_taskID = LockingRRArbiter_4_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_in_0_bits_Typ = LockingRRArbiter_4_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_in_1_valid = LockingRRArbiter_5_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_in_1_bits_RouteID = LockingRRArbiter_5_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_in_1_bits_address = LockingRRArbiter_5_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_in_1_bits_taskID = LockingRRArbiter_5_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_in_1_bits_Typ = LockingRRArbiter_5_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_12_io_out_ready = LockingRRArbiter_16_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_clock = clock;
  assign LockingRRArbiter_13_io_in_0_valid = LockingRRArbiter_6_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_in_0_bits_RouteID = LockingRRArbiter_6_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_in_0_bits_address = LockingRRArbiter_6_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_in_0_bits_taskID = LockingRRArbiter_6_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_in_0_bits_Typ = LockingRRArbiter_6_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_in_1_valid = LockingRRArbiter_7_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_in_1_bits_RouteID = LockingRRArbiter_7_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_in_1_bits_address = LockingRRArbiter_7_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_in_1_bits_taskID = LockingRRArbiter_7_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_in_1_bits_Typ = LockingRRArbiter_7_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_13_io_out_ready = LockingRRArbiter_16_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_clock = clock;
  assign LockingRRArbiter_14_io_in_0_valid = LockingRRArbiter_8_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_in_0_bits_RouteID = LockingRRArbiter_8_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_in_0_bits_address = LockingRRArbiter_8_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_in_0_bits_taskID = LockingRRArbiter_8_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_in_0_bits_Typ = LockingRRArbiter_8_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_in_1_valid = LockingRRArbiter_9_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_in_1_bits_RouteID = LockingRRArbiter_9_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_in_1_bits_address = LockingRRArbiter_9_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_in_1_bits_taskID = LockingRRArbiter_9_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_in_1_bits_Typ = LockingRRArbiter_9_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_14_io_out_ready = LockingRRArbiter_17_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_clock = clock;
  assign LockingRRArbiter_15_io_in_0_valid = LockingRRArbiter_10_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_in_0_bits_RouteID = LockingRRArbiter_10_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_in_0_bits_address = LockingRRArbiter_10_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_in_0_bits_taskID = LockingRRArbiter_10_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_in_0_bits_Typ = LockingRRArbiter_10_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_in_1_valid = LockingRRArbiter_11_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_in_1_bits_RouteID = LockingRRArbiter_11_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_in_1_bits_address = LockingRRArbiter_11_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_in_1_bits_taskID = LockingRRArbiter_11_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_in_1_bits_Typ = LockingRRArbiter_11_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_15_io_out_ready = LockingRRArbiter_18_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_clock = clock;
  assign LockingRRArbiter_16_io_in_0_valid = LockingRRArbiter_12_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_in_0_bits_RouteID = LockingRRArbiter_12_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_in_0_bits_address = LockingRRArbiter_12_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_in_0_bits_taskID = LockingRRArbiter_12_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_in_0_bits_Typ = LockingRRArbiter_12_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_in_1_valid = LockingRRArbiter_13_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_in_1_bits_RouteID = LockingRRArbiter_13_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_in_1_bits_address = LockingRRArbiter_13_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_in_1_bits_taskID = LockingRRArbiter_13_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_in_1_bits_Typ = LockingRRArbiter_13_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_16_io_out_ready = LockingRRArbiter_18_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_17_clock = clock;
  assign LockingRRArbiter_17_io_in_0_valid = LockingRRArbiter_14_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_17_io_in_0_bits_RouteID = LockingRRArbiter_14_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_17_io_in_0_bits_address = LockingRRArbiter_14_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_17_io_in_0_bits_taskID = LockingRRArbiter_14_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_17_io_in_0_bits_Typ = LockingRRArbiter_14_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_17_io_in_1_valid = 1'h0; // @[ArbiterTree.scala 39:67]
  assign LockingRRArbiter_17_io_in_1_bits_RouteID = 16'h0;
  assign LockingRRArbiter_17_io_in_1_bits_address = 32'h0;
  assign LockingRRArbiter_17_io_in_1_bits_taskID = 5'h0;
  assign LockingRRArbiter_17_io_in_1_bits_Typ = 8'h0;
  assign LockingRRArbiter_17_io_out_ready = LockingRRArbiter_19_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_clock = clock;
  assign LockingRRArbiter_18_io_in_0_valid = LockingRRArbiter_15_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_in_0_bits_RouteID = LockingRRArbiter_15_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_in_0_bits_address = LockingRRArbiter_15_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_in_0_bits_taskID = LockingRRArbiter_15_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_in_0_bits_Typ = LockingRRArbiter_15_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_in_1_valid = LockingRRArbiter_16_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_in_1_bits_RouteID = LockingRRArbiter_16_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_in_1_bits_address = LockingRRArbiter_16_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_in_1_bits_taskID = LockingRRArbiter_16_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_in_1_bits_Typ = LockingRRArbiter_16_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_18_io_out_ready = LockingRRArbiter_20_io_in_0_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_19_clock = clock;
  assign LockingRRArbiter_19_io_in_0_valid = LockingRRArbiter_17_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_19_io_in_0_bits_RouteID = LockingRRArbiter_17_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_19_io_in_0_bits_address = LockingRRArbiter_17_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_19_io_in_0_bits_taskID = LockingRRArbiter_17_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_19_io_in_0_bits_Typ = LockingRRArbiter_17_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_19_io_in_1_valid = 1'h0; // @[ArbiterTree.scala 39:67]
  assign LockingRRArbiter_19_io_in_1_bits_RouteID = 16'h0;
  assign LockingRRArbiter_19_io_in_1_bits_address = 32'h0;
  assign LockingRRArbiter_19_io_in_1_bits_taskID = 5'h0;
  assign LockingRRArbiter_19_io_in_1_bits_Typ = 8'h0;
  assign LockingRRArbiter_19_io_out_ready = LockingRRArbiter_20_io_in_1_ready; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_clock = clock;
  assign LockingRRArbiter_20_io_in_0_valid = LockingRRArbiter_18_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_in_0_bits_RouteID = LockingRRArbiter_18_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_in_0_bits_address = LockingRRArbiter_18_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_in_0_bits_taskID = LockingRRArbiter_18_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_in_0_bits_Typ = LockingRRArbiter_18_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_in_1_valid = LockingRRArbiter_19_io_out_valid; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_in_1_bits_RouteID = LockingRRArbiter_19_io_out_bits_RouteID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_in_1_bits_address = LockingRRArbiter_19_io_out_bits_address; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_in_1_bits_taskID = LockingRRArbiter_19_io_out_bits_taskID; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_in_1_bits_Typ = LockingRRArbiter_19_io_out_bits_Typ; // @[ArbiterTree.scala 37:61]
  assign LockingRRArbiter_20_io_out_ready = io_out_ready; // @[ArbiterTree.scala 65:12]
endmodule
module RRArbiter_1(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [15:0] io_in_0_bits_RouteID,
  input  [31:0] io_in_0_bits_data,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [15:0] io_in_1_bits_RouteID,
  input  [31:0] io_in_1_bits_data,
  input         io_out_ready,
  output        io_out_valid,
  output [15:0] io_out_bits_RouteID,
  output [31:0] io_out_bits_data,
  output        io_chosen
);
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Arbiter.scala 67:57]
  wire  _T_5; // @[Arbiter.scala 68:83]
  wire  _T_7; // @[Arbiter.scala 31:68]
  wire  _T_10; // @[Arbiter.scala 31:78]
  wire  _GEN_11; // @[Arbiter.scala 77:27]
  assign _T_3 = 1'h1 > _T_1; // @[Arbiter.scala 67:57]
  assign _T_5 = io_in_1_valid & _T_3; // @[Arbiter.scala 68:83]
  assign _T_7 = _T_5 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_10 = _T_7 == 1'h0; // @[Arbiter.scala 31:78]
  assign _GEN_11 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_5 == 1'h0; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_3 | _T_10; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_RouteID = io_chosen ? io_in_1_bits_RouteID : io_in_0_bits_RouteID; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_5 | _GEN_11; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (io_out_valid) begin
      _T_1 <= io_chosen;
    end
  end
endmodule
module Demux_13(
  input         io_en,
  input  [15:0] io_input_RouteID,
  input  [31:0] io_input_data,
  input         io_sel,
  output        io_outputs_0_valid,
  output [15:0] io_outputs_0_RouteID,
  output [31:0] io_outputs_0_data,
  output        io_outputs_1_valid,
  output [15:0] io_outputs_1_RouteID,
  output [31:0] io_outputs_1_data
);
  wire  _GEN_0; // @[Muxes.scala 29:25]
  assign _GEN_0 = 1'h0 == io_sel; // @[Muxes.scala 29:25]
  assign io_outputs_0_valid = io_en & _GEN_0; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_0_RouteID = io_input_RouteID; // @[Muxes.scala 23:19]
  assign io_outputs_0_data = io_input_data; // @[Muxes.scala 23:19]
  assign io_outputs_1_valid = io_en & io_sel; // @[Muxes.scala 23:19 Muxes.scala 27:27 Muxes.scala 29:25 Muxes.scala 32:27]
  assign io_outputs_1_RouteID = io_input_RouteID; // @[Muxes.scala 23:19]
  assign io_outputs_1_data = io_input_data; // @[Muxes.scala 23:19]
endmodule
module DeMuxTree_1(
  input         clock,
  input         reset,
  output        io_outputs_0_valid,
  output [31:0] io_outputs_0_data,
  output        io_outputs_1_valid,
  output [31:0] io_outputs_1_data,
  output        io_outputs_2_valid,
  output [31:0] io_outputs_2_data,
  output        io_outputs_3_valid,
  output [31:0] io_outputs_3_data,
  output        io_outputs_4_valid,
  output [31:0] io_outputs_4_data,
  output        io_outputs_5_valid,
  output [31:0] io_outputs_5_data,
  output        io_outputs_6_valid,
  output [31:0] io_outputs_6_data,
  output        io_outputs_7_valid,
  output [31:0] io_outputs_7_data,
  output        io_outputs_8_valid,
  output [31:0] io_outputs_8_data,
  output        io_outputs_9_valid,
  output [31:0] io_outputs_9_data,
  output        io_outputs_10_valid,
  output [31:0] io_outputs_10_data,
  output        io_outputs_11_valid,
  output [31:0] io_outputs_11_data,
  output        io_outputs_12_valid,
  output [31:0] io_outputs_12_data,
  output        io_outputs_13_valid,
  output [31:0] io_outputs_13_data,
  output        io_outputs_14_valid,
  output [31:0] io_outputs_14_data,
  output        io_outputs_15_valid,
  output [31:0] io_outputs_15_data,
  output        io_outputs_16_valid,
  output [31:0] io_outputs_16_data,
  output        io_outputs_17_valid,
  output [31:0] io_outputs_17_data,
  output        io_outputs_18_valid,
  output [31:0] io_outputs_18_data,
  input  [15:0] io_input_RouteID,
  input  [31:0] io_input_data,
  input         io_enable
);
  wire  Demux_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_1_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_1_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_1_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_1_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_1_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_1_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_1_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_1_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_1_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_1_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_2_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_2_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_2_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_2_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_2_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_2_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_2_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_2_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_2_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_2_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_3_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_3_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_3_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_3_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_3_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_3_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_3_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_3_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_3_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_3_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_4_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_4_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_4_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_4_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_4_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_4_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_4_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_4_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_4_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_4_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_5_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_5_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_5_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_5_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_5_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_5_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_5_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_5_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_5_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_5_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_6_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_6_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_6_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_6_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_6_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_6_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_6_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_6_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_6_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_6_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_7_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_7_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_7_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_7_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_7_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_7_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_7_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_7_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_7_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_7_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_8_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_8_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_8_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_8_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_8_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_8_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_8_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_8_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_8_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_8_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_9_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_9_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_9_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_9_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_9_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_9_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_9_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_9_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_9_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_9_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_10_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_10_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_10_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_10_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_10_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_10_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_10_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_10_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_10_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_10_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_11_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_11_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_11_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_11_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_11_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_11_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_11_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_11_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_11_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_11_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_12_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_12_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_12_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_12_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_12_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_12_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_12_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_12_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_12_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_12_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_13_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_13_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_13_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_13_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_13_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_13_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_13_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_13_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_13_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_13_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_14_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_14_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_14_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_14_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_14_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_14_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_14_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_14_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_14_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_14_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_15_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_15_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_15_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_15_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_15_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_15_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_15_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_15_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_15_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_15_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_16_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_16_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_16_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_16_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_16_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_16_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_16_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_16_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_16_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_16_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_17_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_17_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_17_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_17_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_17_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_17_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_17_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_17_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_17_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_17_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_18_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_18_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_18_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_18_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_18_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_18_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_18_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_18_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_18_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_18_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_19_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_19_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_19_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_19_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_19_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_19_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_19_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_19_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_19_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_19_io_outputs_1_data; // @[Muxes.scala 91:13]
  wire  Demux_20_io_en; // @[Muxes.scala 91:13]
  wire [15:0] Demux_20_io_input_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_20_io_input_data; // @[Muxes.scala 91:13]
  wire  Demux_20_io_sel; // @[Muxes.scala 91:13]
  wire  Demux_20_io_outputs_0_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_20_io_outputs_0_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_20_io_outputs_0_data; // @[Muxes.scala 91:13]
  wire  Demux_20_io_outputs_1_valid; // @[Muxes.scala 91:13]
  wire [15:0] Demux_20_io_outputs_1_RouteID; // @[Muxes.scala 91:13]
  wire [31:0] Demux_20_io_outputs_1_data; // @[Muxes.scala 91:13]
  reg [15:0] _T_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_0;
  reg [31:0] _T_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_1;
  reg  _T_1; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_2;
  reg [15:0] _T_3_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_3;
  reg [31:0] _T_3_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_4;
  reg  _T_4; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_5;
  reg [15:0] _T_6_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_6;
  reg [31:0] _T_6_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_7;
  reg  _T_7; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_8;
  reg [15:0] _T_9_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_9;
  reg [31:0] _T_9_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_10;
  reg  _T_10; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_11;
  reg [15:0] _T_12_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_12;
  reg [31:0] _T_12_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_13;
  reg  _T_13; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_14;
  reg [15:0] _T_15_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_15;
  reg [31:0] _T_15_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_16;
  reg  _T_16; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_17;
  reg [15:0] _T_18_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_18;
  reg [31:0] _T_18_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_19;
  reg  _T_19; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_20;
  reg [15:0] _T_21_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_21;
  reg [31:0] _T_21_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_22;
  reg  _T_22; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_23;
  reg [15:0] _T_24_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_24;
  reg [31:0] _T_24_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_25;
  reg  _T_25; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_26;
  reg [15:0] _T_27_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_27;
  reg [31:0] _T_27_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_28;
  reg  _T_28; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_29;
  reg [15:0] _T_30_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_30;
  reg [31:0] _T_30_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_31;
  reg  _T_31; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_32;
  reg [15:0] _T_33_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_33;
  reg [31:0] _T_33_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_34;
  reg  _T_34; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_35;
  reg [15:0] _T_36_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_36;
  reg [31:0] _T_36_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_37;
  reg  _T_37; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_38;
  reg [15:0] _T_39_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_39;
  reg [31:0] _T_39_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_40;
  reg  _T_40; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_41;
  reg [15:0] _T_42_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_42;
  reg [31:0] _T_42_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_43;
  reg  _T_43; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_44;
  reg [15:0] _T_45_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_45;
  reg [31:0] _T_45_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_46;
  reg  _T_46; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_47;
  reg [15:0] _T_48_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_48;
  reg [31:0] _T_48_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_49;
  reg  _T_49; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_50;
  reg [15:0] _T_51_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_51;
  reg [31:0] _T_51_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_52;
  reg  _T_52; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_53;
  reg [15:0] _T_54_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_54;
  reg [31:0] _T_54_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_55;
  reg  _T_55; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_56;
  reg [15:0] _T_57_RouteID; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_57;
  reg [31:0] _T_57_data; // @[Muxes.scala 102:36]
  reg [31:0] _RAND_58;
  reg  _T_58; // @[Muxes.scala 103:36]
  reg [31:0] _RAND_59;
  Demux_13 Demux ( // @[Muxes.scala 91:13]
    .io_en(Demux_io_en),
    .io_input_RouteID(Demux_io_input_RouteID),
    .io_input_data(Demux_io_input_data),
    .io_sel(Demux_io_sel),
    .io_outputs_0_valid(Demux_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_io_outputs_0_data),
    .io_outputs_1_valid(Demux_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_io_outputs_1_data)
  );
  Demux_13 Demux_1 ( // @[Muxes.scala 91:13]
    .io_en(Demux_1_io_en),
    .io_input_RouteID(Demux_1_io_input_RouteID),
    .io_input_data(Demux_1_io_input_data),
    .io_sel(Demux_1_io_sel),
    .io_outputs_0_valid(Demux_1_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_1_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_1_io_outputs_0_data),
    .io_outputs_1_valid(Demux_1_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_1_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_1_io_outputs_1_data)
  );
  Demux_13 Demux_2 ( // @[Muxes.scala 91:13]
    .io_en(Demux_2_io_en),
    .io_input_RouteID(Demux_2_io_input_RouteID),
    .io_input_data(Demux_2_io_input_data),
    .io_sel(Demux_2_io_sel),
    .io_outputs_0_valid(Demux_2_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_2_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_2_io_outputs_0_data),
    .io_outputs_1_valid(Demux_2_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_2_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_2_io_outputs_1_data)
  );
  Demux_13 Demux_3 ( // @[Muxes.scala 91:13]
    .io_en(Demux_3_io_en),
    .io_input_RouteID(Demux_3_io_input_RouteID),
    .io_input_data(Demux_3_io_input_data),
    .io_sel(Demux_3_io_sel),
    .io_outputs_0_valid(Demux_3_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_3_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_3_io_outputs_0_data),
    .io_outputs_1_valid(Demux_3_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_3_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_3_io_outputs_1_data)
  );
  Demux_13 Demux_4 ( // @[Muxes.scala 91:13]
    .io_en(Demux_4_io_en),
    .io_input_RouteID(Demux_4_io_input_RouteID),
    .io_input_data(Demux_4_io_input_data),
    .io_sel(Demux_4_io_sel),
    .io_outputs_0_valid(Demux_4_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_4_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_4_io_outputs_0_data),
    .io_outputs_1_valid(Demux_4_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_4_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_4_io_outputs_1_data)
  );
  Demux_13 Demux_5 ( // @[Muxes.scala 91:13]
    .io_en(Demux_5_io_en),
    .io_input_RouteID(Demux_5_io_input_RouteID),
    .io_input_data(Demux_5_io_input_data),
    .io_sel(Demux_5_io_sel),
    .io_outputs_0_valid(Demux_5_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_5_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_5_io_outputs_0_data),
    .io_outputs_1_valid(Demux_5_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_5_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_5_io_outputs_1_data)
  );
  Demux_13 Demux_6 ( // @[Muxes.scala 91:13]
    .io_en(Demux_6_io_en),
    .io_input_RouteID(Demux_6_io_input_RouteID),
    .io_input_data(Demux_6_io_input_data),
    .io_sel(Demux_6_io_sel),
    .io_outputs_0_valid(Demux_6_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_6_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_6_io_outputs_0_data),
    .io_outputs_1_valid(Demux_6_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_6_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_6_io_outputs_1_data)
  );
  Demux_13 Demux_7 ( // @[Muxes.scala 91:13]
    .io_en(Demux_7_io_en),
    .io_input_RouteID(Demux_7_io_input_RouteID),
    .io_input_data(Demux_7_io_input_data),
    .io_sel(Demux_7_io_sel),
    .io_outputs_0_valid(Demux_7_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_7_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_7_io_outputs_0_data),
    .io_outputs_1_valid(Demux_7_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_7_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_7_io_outputs_1_data)
  );
  Demux_13 Demux_8 ( // @[Muxes.scala 91:13]
    .io_en(Demux_8_io_en),
    .io_input_RouteID(Demux_8_io_input_RouteID),
    .io_input_data(Demux_8_io_input_data),
    .io_sel(Demux_8_io_sel),
    .io_outputs_0_valid(Demux_8_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_8_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_8_io_outputs_0_data),
    .io_outputs_1_valid(Demux_8_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_8_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_8_io_outputs_1_data)
  );
  Demux_13 Demux_9 ( // @[Muxes.scala 91:13]
    .io_en(Demux_9_io_en),
    .io_input_RouteID(Demux_9_io_input_RouteID),
    .io_input_data(Demux_9_io_input_data),
    .io_sel(Demux_9_io_sel),
    .io_outputs_0_valid(Demux_9_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_9_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_9_io_outputs_0_data),
    .io_outputs_1_valid(Demux_9_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_9_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_9_io_outputs_1_data)
  );
  Demux_13 Demux_10 ( // @[Muxes.scala 91:13]
    .io_en(Demux_10_io_en),
    .io_input_RouteID(Demux_10_io_input_RouteID),
    .io_input_data(Demux_10_io_input_data),
    .io_sel(Demux_10_io_sel),
    .io_outputs_0_valid(Demux_10_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_10_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_10_io_outputs_0_data),
    .io_outputs_1_valid(Demux_10_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_10_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_10_io_outputs_1_data)
  );
  Demux_13 Demux_11 ( // @[Muxes.scala 91:13]
    .io_en(Demux_11_io_en),
    .io_input_RouteID(Demux_11_io_input_RouteID),
    .io_input_data(Demux_11_io_input_data),
    .io_sel(Demux_11_io_sel),
    .io_outputs_0_valid(Demux_11_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_11_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_11_io_outputs_0_data),
    .io_outputs_1_valid(Demux_11_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_11_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_11_io_outputs_1_data)
  );
  Demux_13 Demux_12 ( // @[Muxes.scala 91:13]
    .io_en(Demux_12_io_en),
    .io_input_RouteID(Demux_12_io_input_RouteID),
    .io_input_data(Demux_12_io_input_data),
    .io_sel(Demux_12_io_sel),
    .io_outputs_0_valid(Demux_12_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_12_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_12_io_outputs_0_data),
    .io_outputs_1_valid(Demux_12_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_12_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_12_io_outputs_1_data)
  );
  Demux_13 Demux_13 ( // @[Muxes.scala 91:13]
    .io_en(Demux_13_io_en),
    .io_input_RouteID(Demux_13_io_input_RouteID),
    .io_input_data(Demux_13_io_input_data),
    .io_sel(Demux_13_io_sel),
    .io_outputs_0_valid(Demux_13_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_13_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_13_io_outputs_0_data),
    .io_outputs_1_valid(Demux_13_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_13_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_13_io_outputs_1_data)
  );
  Demux_13 Demux_14 ( // @[Muxes.scala 91:13]
    .io_en(Demux_14_io_en),
    .io_input_RouteID(Demux_14_io_input_RouteID),
    .io_input_data(Demux_14_io_input_data),
    .io_sel(Demux_14_io_sel),
    .io_outputs_0_valid(Demux_14_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_14_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_14_io_outputs_0_data),
    .io_outputs_1_valid(Demux_14_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_14_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_14_io_outputs_1_data)
  );
  Demux_13 Demux_15 ( // @[Muxes.scala 91:13]
    .io_en(Demux_15_io_en),
    .io_input_RouteID(Demux_15_io_input_RouteID),
    .io_input_data(Demux_15_io_input_data),
    .io_sel(Demux_15_io_sel),
    .io_outputs_0_valid(Demux_15_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_15_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_15_io_outputs_0_data),
    .io_outputs_1_valid(Demux_15_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_15_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_15_io_outputs_1_data)
  );
  Demux_13 Demux_16 ( // @[Muxes.scala 91:13]
    .io_en(Demux_16_io_en),
    .io_input_RouteID(Demux_16_io_input_RouteID),
    .io_input_data(Demux_16_io_input_data),
    .io_sel(Demux_16_io_sel),
    .io_outputs_0_valid(Demux_16_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_16_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_16_io_outputs_0_data),
    .io_outputs_1_valid(Demux_16_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_16_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_16_io_outputs_1_data)
  );
  Demux_13 Demux_17 ( // @[Muxes.scala 91:13]
    .io_en(Demux_17_io_en),
    .io_input_RouteID(Demux_17_io_input_RouteID),
    .io_input_data(Demux_17_io_input_data),
    .io_sel(Demux_17_io_sel),
    .io_outputs_0_valid(Demux_17_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_17_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_17_io_outputs_0_data),
    .io_outputs_1_valid(Demux_17_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_17_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_17_io_outputs_1_data)
  );
  Demux_13 Demux_18 ( // @[Muxes.scala 91:13]
    .io_en(Demux_18_io_en),
    .io_input_RouteID(Demux_18_io_input_RouteID),
    .io_input_data(Demux_18_io_input_data),
    .io_sel(Demux_18_io_sel),
    .io_outputs_0_valid(Demux_18_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_18_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_18_io_outputs_0_data),
    .io_outputs_1_valid(Demux_18_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_18_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_18_io_outputs_1_data)
  );
  Demux_13 Demux_19 ( // @[Muxes.scala 91:13]
    .io_en(Demux_19_io_en),
    .io_input_RouteID(Demux_19_io_input_RouteID),
    .io_input_data(Demux_19_io_input_data),
    .io_sel(Demux_19_io_sel),
    .io_outputs_0_valid(Demux_19_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_19_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_19_io_outputs_0_data),
    .io_outputs_1_valid(Demux_19_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_19_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_19_io_outputs_1_data)
  );
  Demux_13 Demux_20 ( // @[Muxes.scala 91:13]
    .io_en(Demux_20_io_en),
    .io_input_RouteID(Demux_20_io_input_RouteID),
    .io_input_data(Demux_20_io_input_data),
    .io_sel(Demux_20_io_sel),
    .io_outputs_0_valid(Demux_20_io_outputs_0_valid),
    .io_outputs_0_RouteID(Demux_20_io_outputs_0_RouteID),
    .io_outputs_0_data(Demux_20_io_outputs_0_data),
    .io_outputs_1_valid(Demux_20_io_outputs_1_valid),
    .io_outputs_1_RouteID(Demux_20_io_outputs_1_RouteID),
    .io_outputs_1_data(Demux_20_io_outputs_1_data)
  );
  assign io_outputs_0_valid = Demux_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_0_data = Demux_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_1_valid = Demux_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_1_data = Demux_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_2_valid = Demux_1_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_2_data = Demux_1_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_3_valid = Demux_1_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_3_data = Demux_1_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_4_valid = Demux_2_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_4_data = Demux_2_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_5_valid = Demux_2_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_5_data = Demux_2_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_6_valid = Demux_3_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_6_data = Demux_3_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_7_valid = Demux_3_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_7_data = Demux_3_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_8_valid = Demux_4_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_8_data = Demux_4_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_9_valid = Demux_4_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_9_data = Demux_4_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_10_valid = Demux_5_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_10_data = Demux_5_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_11_valid = Demux_5_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_11_data = Demux_5_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_12_valid = Demux_6_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_12_data = Demux_6_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_13_valid = Demux_6_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_13_data = Demux_6_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_14_valid = Demux_7_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_14_data = Demux_7_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_15_valid = Demux_7_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_15_data = Demux_7_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_16_valid = Demux_8_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_16_data = Demux_8_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign io_outputs_17_valid = Demux_8_io_outputs_1_valid; // @[Muxes.scala 119:25]
  assign io_outputs_17_data = Demux_8_io_outputs_1_data; // @[Muxes.scala 119:25]
  assign io_outputs_18_valid = Demux_9_io_outputs_0_valid; // @[Muxes.scala 119:25]
  assign io_outputs_18_data = Demux_9_io_outputs_0_data; // @[Muxes.scala 119:25]
  assign Demux_io_en = _T_1; // @[Muxes.scala 105:20]
  assign Demux_io_input_RouteID = _T_RouteID; // @[Muxes.scala 104:23]
  assign Demux_io_input_data = _T_data; // @[Muxes.scala 104:23]
  assign Demux_io_sel = _T_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_1_io_en = _T_4; // @[Muxes.scala 105:20]
  assign Demux_1_io_input_RouteID = _T_3_RouteID; // @[Muxes.scala 104:23]
  assign Demux_1_io_input_data = _T_3_data; // @[Muxes.scala 104:23]
  assign Demux_1_io_sel = _T_3_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_2_io_en = _T_7; // @[Muxes.scala 105:20]
  assign Demux_2_io_input_RouteID = _T_6_RouteID; // @[Muxes.scala 104:23]
  assign Demux_2_io_input_data = _T_6_data; // @[Muxes.scala 104:23]
  assign Demux_2_io_sel = _T_6_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_3_io_en = _T_10; // @[Muxes.scala 105:20]
  assign Demux_3_io_input_RouteID = _T_9_RouteID; // @[Muxes.scala 104:23]
  assign Demux_3_io_input_data = _T_9_data; // @[Muxes.scala 104:23]
  assign Demux_3_io_sel = _T_9_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_4_io_en = _T_13; // @[Muxes.scala 105:20]
  assign Demux_4_io_input_RouteID = _T_12_RouteID; // @[Muxes.scala 104:23]
  assign Demux_4_io_input_data = _T_12_data; // @[Muxes.scala 104:23]
  assign Demux_4_io_sel = _T_12_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_5_io_en = _T_16; // @[Muxes.scala 105:20]
  assign Demux_5_io_input_RouteID = _T_15_RouteID; // @[Muxes.scala 104:23]
  assign Demux_5_io_input_data = _T_15_data; // @[Muxes.scala 104:23]
  assign Demux_5_io_sel = _T_15_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_6_io_en = _T_19; // @[Muxes.scala 105:20]
  assign Demux_6_io_input_RouteID = _T_18_RouteID; // @[Muxes.scala 104:23]
  assign Demux_6_io_input_data = _T_18_data; // @[Muxes.scala 104:23]
  assign Demux_6_io_sel = _T_18_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_7_io_en = _T_22; // @[Muxes.scala 105:20]
  assign Demux_7_io_input_RouteID = _T_21_RouteID; // @[Muxes.scala 104:23]
  assign Demux_7_io_input_data = _T_21_data; // @[Muxes.scala 104:23]
  assign Demux_7_io_sel = _T_21_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_8_io_en = _T_25; // @[Muxes.scala 105:20]
  assign Demux_8_io_input_RouteID = _T_24_RouteID; // @[Muxes.scala 104:23]
  assign Demux_8_io_input_data = _T_24_data; // @[Muxes.scala 104:23]
  assign Demux_8_io_sel = _T_24_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_9_io_en = _T_28; // @[Muxes.scala 105:20]
  assign Demux_9_io_input_RouteID = _T_27_RouteID; // @[Muxes.scala 104:23]
  assign Demux_9_io_input_data = _T_27_data; // @[Muxes.scala 104:23]
  assign Demux_9_io_sel = _T_27_RouteID[0]; // @[Muxes.scala 106:21]
  assign Demux_10_io_en = _T_31; // @[Muxes.scala 105:20]
  assign Demux_10_io_input_RouteID = _T_30_RouteID; // @[Muxes.scala 104:23]
  assign Demux_10_io_input_data = _T_30_data; // @[Muxes.scala 104:23]
  assign Demux_10_io_sel = _T_30_RouteID[1]; // @[Muxes.scala 106:21]
  assign Demux_11_io_en = _T_34; // @[Muxes.scala 105:20]
  assign Demux_11_io_input_RouteID = _T_33_RouteID; // @[Muxes.scala 104:23]
  assign Demux_11_io_input_data = _T_33_data; // @[Muxes.scala 104:23]
  assign Demux_11_io_sel = _T_33_RouteID[1]; // @[Muxes.scala 106:21]
  assign Demux_12_io_en = _T_37; // @[Muxes.scala 105:20]
  assign Demux_12_io_input_RouteID = _T_36_RouteID; // @[Muxes.scala 104:23]
  assign Demux_12_io_input_data = _T_36_data; // @[Muxes.scala 104:23]
  assign Demux_12_io_sel = _T_36_RouteID[1]; // @[Muxes.scala 106:21]
  assign Demux_13_io_en = _T_40; // @[Muxes.scala 105:20]
  assign Demux_13_io_input_RouteID = _T_39_RouteID; // @[Muxes.scala 104:23]
  assign Demux_13_io_input_data = _T_39_data; // @[Muxes.scala 104:23]
  assign Demux_13_io_sel = _T_39_RouteID[1]; // @[Muxes.scala 106:21]
  assign Demux_14_io_en = _T_43; // @[Muxes.scala 105:20]
  assign Demux_14_io_input_RouteID = _T_42_RouteID; // @[Muxes.scala 104:23]
  assign Demux_14_io_input_data = _T_42_data; // @[Muxes.scala 104:23]
  assign Demux_14_io_sel = _T_42_RouteID[1]; // @[Muxes.scala 106:21]
  assign Demux_15_io_en = _T_46; // @[Muxes.scala 105:20]
  assign Demux_15_io_input_RouteID = _T_45_RouteID; // @[Muxes.scala 104:23]
  assign Demux_15_io_input_data = _T_45_data; // @[Muxes.scala 104:23]
  assign Demux_15_io_sel = _T_45_RouteID[2]; // @[Muxes.scala 106:21]
  assign Demux_16_io_en = _T_49; // @[Muxes.scala 105:20]
  assign Demux_16_io_input_RouteID = _T_48_RouteID; // @[Muxes.scala 104:23]
  assign Demux_16_io_input_data = _T_48_data; // @[Muxes.scala 104:23]
  assign Demux_16_io_sel = _T_48_RouteID[2]; // @[Muxes.scala 106:21]
  assign Demux_17_io_en = _T_52; // @[Muxes.scala 105:20]
  assign Demux_17_io_input_RouteID = _T_51_RouteID; // @[Muxes.scala 104:23]
  assign Demux_17_io_input_data = _T_51_data; // @[Muxes.scala 104:23]
  assign Demux_17_io_sel = _T_51_RouteID[2]; // @[Muxes.scala 106:21]
  assign Demux_18_io_en = _T_55; // @[Muxes.scala 105:20]
  assign Demux_18_io_input_RouteID = _T_54_RouteID; // @[Muxes.scala 104:23]
  assign Demux_18_io_input_data = _T_54_data; // @[Muxes.scala 104:23]
  assign Demux_18_io_sel = _T_54_RouteID[3]; // @[Muxes.scala 106:21]
  assign Demux_19_io_en = _T_58; // @[Muxes.scala 105:20]
  assign Demux_19_io_input_RouteID = _T_57_RouteID; // @[Muxes.scala 104:23]
  assign Demux_19_io_input_data = _T_57_data; // @[Muxes.scala 104:23]
  assign Demux_19_io_sel = _T_57_RouteID[3]; // @[Muxes.scala 106:21]
  assign Demux_20_io_en = io_enable; // @[Muxes.scala 135:14]
  assign Demux_20_io_input_RouteID = io_input_RouteID; // @[Muxes.scala 134:17]
  assign Demux_20_io_input_data = io_input_data; // @[Muxes.scala 134:17]
  assign Demux_20_io_sel = io_input_RouteID[4]; // @[Muxes.scala 136:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_RouteID = _RAND_0[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_3_RouteID = _RAND_3[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_3_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_4 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_6_RouteID = _RAND_6[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_6_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_7 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_9_RouteID = _RAND_9[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_9_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_10 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_12_RouteID = _RAND_12[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_12_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_13 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T_15_RouteID = _RAND_15[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_15_data = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_16 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_18_RouteID = _RAND_18[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  _T_18_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_19 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_21_RouteID = _RAND_21[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_21_data = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_22 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_24_RouteID = _RAND_24[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_24_data = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_25 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_27_RouteID = _RAND_27[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_27_data = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_28 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_30_RouteID = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_30_data = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_31 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_33_RouteID = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_33_data = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_34 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_36_RouteID = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_36_data = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_37 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_39_RouteID = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_39_data = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_40 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_42_RouteID = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_42_data = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_43 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_45_RouteID = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_45_data = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_46 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_48_RouteID = _RAND_48[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_48_data = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_49 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_51_RouteID = _RAND_51[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_51_data = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_52 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_54_RouteID = _RAND_54[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_54_data = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_55 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_57_RouteID = _RAND_57[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_57_data = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_58 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    _T_RouteID <= Demux_10_io_outputs_0_RouteID;
    _T_data <= Demux_10_io_outputs_0_data;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= Demux_10_io_outputs_0_valid;
    end
    _T_3_RouteID <= Demux_10_io_outputs_1_RouteID;
    _T_3_data <= Demux_10_io_outputs_1_data;
    if (reset) begin
      _T_4 <= 1'h0;
    end else begin
      _T_4 <= Demux_10_io_outputs_1_valid;
    end
    _T_6_RouteID <= Demux_11_io_outputs_0_RouteID;
    _T_6_data <= Demux_11_io_outputs_0_data;
    if (reset) begin
      _T_7 <= 1'h0;
    end else begin
      _T_7 <= Demux_11_io_outputs_0_valid;
    end
    _T_9_RouteID <= Demux_11_io_outputs_1_RouteID;
    _T_9_data <= Demux_11_io_outputs_1_data;
    if (reset) begin
      _T_10 <= 1'h0;
    end else begin
      _T_10 <= Demux_11_io_outputs_1_valid;
    end
    _T_12_RouteID <= Demux_12_io_outputs_0_RouteID;
    _T_12_data <= Demux_12_io_outputs_0_data;
    if (reset) begin
      _T_13 <= 1'h0;
    end else begin
      _T_13 <= Demux_12_io_outputs_0_valid;
    end
    _T_15_RouteID <= Demux_12_io_outputs_1_RouteID;
    _T_15_data <= Demux_12_io_outputs_1_data;
    if (reset) begin
      _T_16 <= 1'h0;
    end else begin
      _T_16 <= Demux_12_io_outputs_1_valid;
    end
    _T_18_RouteID <= Demux_13_io_outputs_0_RouteID;
    _T_18_data <= Demux_13_io_outputs_0_data;
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      _T_19 <= Demux_13_io_outputs_0_valid;
    end
    _T_21_RouteID <= Demux_13_io_outputs_1_RouteID;
    _T_21_data <= Demux_13_io_outputs_1_data;
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      _T_22 <= Demux_13_io_outputs_1_valid;
    end
    _T_24_RouteID <= Demux_14_io_outputs_0_RouteID;
    _T_24_data <= Demux_14_io_outputs_0_data;
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      _T_25 <= Demux_14_io_outputs_0_valid;
    end
    _T_27_RouteID <= Demux_14_io_outputs_1_RouteID;
    _T_27_data <= Demux_14_io_outputs_1_data;
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      _T_28 <= Demux_14_io_outputs_1_valid;
    end
    _T_30_RouteID <= Demux_15_io_outputs_0_RouteID;
    _T_30_data <= Demux_15_io_outputs_0_data;
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      _T_31 <= Demux_15_io_outputs_0_valid;
    end
    _T_33_RouteID <= Demux_15_io_outputs_1_RouteID;
    _T_33_data <= Demux_15_io_outputs_1_data;
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      _T_34 <= Demux_15_io_outputs_1_valid;
    end
    _T_36_RouteID <= Demux_16_io_outputs_0_RouteID;
    _T_36_data <= Demux_16_io_outputs_0_data;
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      _T_37 <= Demux_16_io_outputs_0_valid;
    end
    _T_39_RouteID <= Demux_16_io_outputs_1_RouteID;
    _T_39_data <= Demux_16_io_outputs_1_data;
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      _T_40 <= Demux_16_io_outputs_1_valid;
    end
    _T_42_RouteID <= Demux_17_io_outputs_0_RouteID;
    _T_42_data <= Demux_17_io_outputs_0_data;
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      _T_43 <= Demux_17_io_outputs_0_valid;
    end
    _T_45_RouteID <= Demux_18_io_outputs_0_RouteID;
    _T_45_data <= Demux_18_io_outputs_0_data;
    if (reset) begin
      _T_46 <= 1'h0;
    end else begin
      _T_46 <= Demux_18_io_outputs_0_valid;
    end
    _T_48_RouteID <= Demux_18_io_outputs_1_RouteID;
    _T_48_data <= Demux_18_io_outputs_1_data;
    if (reset) begin
      _T_49 <= 1'h0;
    end else begin
      _T_49 <= Demux_18_io_outputs_1_valid;
    end
    _T_51_RouteID <= Demux_19_io_outputs_0_RouteID;
    _T_51_data <= Demux_19_io_outputs_0_data;
    if (reset) begin
      _T_52 <= 1'h0;
    end else begin
      _T_52 <= Demux_19_io_outputs_0_valid;
    end
    _T_54_RouteID <= Demux_20_io_outputs_0_RouteID;
    _T_54_data <= Demux_20_io_outputs_0_data;
    if (reset) begin
      _T_55 <= 1'h0;
    end else begin
      _T_55 <= Demux_20_io_outputs_0_valid;
    end
    _T_57_RouteID <= Demux_20_io_outputs_1_RouteID;
    _T_57_data <= Demux_20_io_outputs_1_data;
    if (reset) begin
      _T_58 <= 1'h0;
    end else begin
      _T_58 <= Demux_20_io_outputs_1_valid;
    end
  end
endmodule
module ReadTableEntry(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [15:0] io_NodeReq_bits_RouteID,
  input  [31:0] io_NodeReq_bits_address,
  input  [4:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_data,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output [31:0] io_output_bits_data,
  output        io_free
);
  reg  ID; // @[ReadMemoryController.scala 49:19]
  reg [31:0] _RAND_0;
  reg [15:0] request_R_RouteID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_1;
  reg [31:0] request_R_address; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_2;
  reg [4:0] request_R_taskID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_3;
  reg [7:0] request_R_Typ; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_4;
  reg [63:0] bitmask; // @[ReadMemoryController.scala 56:29]
  reg [63:0] _RAND_5;
  reg [7:0] sendbytemask; // @[ReadMemoryController.scala 58:29]
  reg [31:0] _RAND_6;
  reg [31:0] ReqAddress; // @[ReadMemoryController.scala 62:27]
  reg [31:0] _RAND_7;
  reg  ptr; // @[ReadMemoryController.scala 66:27]
  reg [31:0] _RAND_8;
  reg [31:0] linebuffer_0; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_9;
  reg [31:0] linebuffer_1; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[ReadMemoryController.scala 73:68]
  reg [31:0] _RAND_11;
  wire [2:0] _T_6; // @[Cat.scala 29:58]
  wire [31:0] _GEN_57; // @[ReadMemoryController.scala 96:37]
  reg  isWrite; // @[ReadMemoryController.scala 100:24]
  reg [31:0] _RAND_12;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire [29:0] _T_10; // @[ReadMemoryController.scala 115:44]
  wire [31:0] _T_11; // @[ReadMemoryController.scala 115:69]
  wire  _T_12; // @[helpers.scala 27:24]
  wire  _T_13; // @[helpers.scala 27:47]
  wire  _T_14; // @[helpers.scala 27:40]
  wire  _T_16; // @[helpers.scala 28:15]
  wire  _T_17; // @[helpers.scala 28:38]
  wire  _T_18; // @[helpers.scala 28:31]
  wire  _T_20; // @[helpers.scala 29:17]
  wire  _T_21; // @[helpers.scala 29:40]
  wire  _T_22; // @[helpers.scala 29:33]
  wire [63:0] _T_25; // @[helpers.scala 29:12]
  wire [63:0] _T_26; // @[helpers.scala 28:10]
  wire [63:0] _T_27; // @[helpers.scala 27:19]
  wire [1:0] _T_28; // @[helpers.scala 39:32]
  wire [4:0] _T_29; // @[Cat.scala 29:58]
  wire [94:0] _GEN_58; // @[helpers.scala 40:26]
  wire [94:0] _T_30; // @[helpers.scala 40:26]
  wire [7:0] _T_43; // @[helpers.scala 50:12]
  wire [7:0] _T_44; // @[helpers.scala 49:10]
  wire [7:0] _T_45; // @[helpers.scala 48:19]
  wire [10:0] _GEN_59; // @[helpers.scala 20:26]
  wire [10:0] _T_47; // @[helpers.scala 20:26]
  wire [94:0] _GEN_5; // @[ReadMemoryController.scala 111:28]
  wire [10:0] _GEN_6; // @[ReadMemoryController.scala 111:28]
  wire  _T_48; // @[Conditional.scala 37:30]
  wire  _T_50; // @[Conditional.scala 37:30]
  wire [3:0] _T_51; // @[ReadMemoryController.scala 144:38]
  wire [10:0] _GEN_8; // @[ReadMemoryController.scala 142:29]
  wire  _T_52; // @[Conditional.scala 37:30]
  wire  _T_54; // @[ReadMemoryController.scala 154:20]
  wire  _T_55; // @[ReadMemoryController.scala 156:27]
  wire  _T_56; // @[Conditional.scala 37:30]
  wire [63:0] _T_57; // @[ReadMemoryController.scala 165:29]
  wire [63:0] _T_58; // @[ReadMemoryController.scala 165:36]
  wire [1:0] _T_59; // @[ReadMemoryController.scala 165:71]
  wire [4:0] _T_60; // @[Cat.scala 29:58]
  wire [63:0] _T_61; // @[ReadMemoryController.scala 165:47]
  wire  _T_62; // @[helpers.scala 63:30]
  wire [63:0] _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_31; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_42; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_53; // @[Conditional.scala 40:58]
  wire [31:0] output_; // @[ReadMemoryController.scala 165:14]
  wire  _T_63; // @[helpers.scala 63:57]
  wire [15:0] _T_65; // @[Bitwise.scala 71:12]
  wire [15:0] _T_66; // @[helpers.scala 63:68]
  wire [31:0] _T_67; // @[Cat.scala 29:58]
  wire  _T_68; // @[helpers.scala 64:22]
  wire [31:0] _T_71; // @[Cat.scala 29:58]
  wire  _T_72; // @[helpers.scala 65:24]
  wire  _T_73; // @[helpers.scala 65:51]
  wire [23:0] _T_75; // @[Bitwise.scala 71:12]
  wire [7:0] _T_76; // @[helpers.scala 65:61]
  wire [31:0] _T_77; // @[Cat.scala 29:58]
  wire  _T_78; // @[helpers.scala 66:26]
  wire [31:0] _T_81; // @[Cat.scala 29:58]
  wire [31:0] _T_83; // @[helpers.scala 66:14]
  wire [31:0] _T_84; // @[helpers.scala 65:12]
  wire [31:0] _T_85; // @[helpers.scala 64:10]
  wire [31:0] _T_86; // @[helpers.scala 63:18]
  wire [31:0] _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_43; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_48; // @[Conditional.scala 40:58]
  assign _T_6 = {ptr,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_57 = {{29'd0}, _T_6}; // @[ReadMemoryController.scala 96:37]
  assign _T_9 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_NodeReq_bits_address[31:2]; // @[ReadMemoryController.scala 115:44]
  assign _T_11 = {_T_10, 2'h0}; // @[ReadMemoryController.scala 115:69]
  assign _T_12 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_13 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_14 = _T_12 | _T_13; // @[helpers.scala 27:40]
  assign _T_16 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_17 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_18 = _T_16 | _T_17; // @[helpers.scala 28:31]
  assign _T_20 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_21 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_22 = _T_20 | _T_21; // @[helpers.scala 29:33]
  assign _T_25 = _T_22 ? 64'hffffffff : 64'hffffffffffffffff; // @[helpers.scala 29:12]
  assign _T_26 = _T_18 ? 64'hff : _T_25; // @[helpers.scala 28:10]
  assign _T_27 = _T_14 ? 64'hffff : _T_26; // @[helpers.scala 27:19]
  assign _T_28 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_29 = {_T_28,3'h0}; // @[Cat.scala 29:58]
  assign _GEN_58 = {{31'd0}, _T_27}; // @[helpers.scala 40:26]
  assign _T_30 = _GEN_58 << _T_29; // @[helpers.scala 40:26]
  assign _T_43 = _T_22 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_44 = _T_18 ? 8'h1 : _T_43; // @[helpers.scala 49:10]
  assign _T_45 = _T_14 ? 8'h3 : _T_44; // @[helpers.scala 48:19]
  assign _GEN_59 = {{3'd0}, _T_45}; // @[helpers.scala 20:26]
  assign _T_47 = _GEN_59 << _T_28; // @[helpers.scala 20:26]
  assign _GEN_5 = _T_9 ? _T_30 : {{31'd0}, bitmask}; // @[ReadMemoryController.scala 111:28]
  assign _GEN_6 = _T_9 ? _T_47 : {{3'd0}, sendbytemask}; // @[ReadMemoryController.scala 111:28]
  assign _T_48 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_50 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_51 = sendbytemask[7:4]; // @[ReadMemoryController.scala 144:38]
  assign _GEN_8 = io_MemReq_ready ? {{7'd0}, _T_51} : _GEN_6; // @[ReadMemoryController.scala 142:29]
  assign _T_52 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_54 = ptr + 1'h1; // @[ReadMemoryController.scala 154:20]
  assign _T_55 = sendbytemask == 8'h0; // @[ReadMemoryController.scala 156:27]
  assign _T_56 = 2'h3 == state; // @[Conditional.scala 37:30]
  assign _T_57 = {linebuffer_1,linebuffer_0}; // @[ReadMemoryController.scala 165:29]
  assign _T_58 = _T_57 & bitmask; // @[ReadMemoryController.scala 165:36]
  assign _T_59 = request_R_address[1:0]; // @[ReadMemoryController.scala 165:71]
  assign _T_60 = {_T_59,3'h0}; // @[Cat.scala 29:58]
  assign _T_61 = _T_58 >> _T_60; // @[ReadMemoryController.scala 165:47]
  assign _T_62 = request_R_Typ == 8'h2; // @[helpers.scala 63:30]
  assign _GEN_20 = _T_56 ? _T_61 : 64'h0; // @[Conditional.scala 39:67]
  assign _GEN_31 = _T_52 ? 64'h0 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_50 ? 64'h0 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_53 = _T_48 ? 64'h0 : _GEN_42; // @[Conditional.scala 40:58]
  assign output_ = _GEN_53[31:0]; // @[ReadMemoryController.scala 165:14]
  assign _T_63 = output_[15]; // @[helpers.scala 63:57]
  assign _T_65 = _T_63 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_66 = output_[15:0]; // @[helpers.scala 63:68]
  assign _T_67 = {_T_65,_T_66}; // @[Cat.scala 29:58]
  assign _T_68 = request_R_Typ == 8'h6; // @[helpers.scala 64:22]
  assign _T_71 = {16'h0,_T_66}; // @[Cat.scala 29:58]
  assign _T_72 = request_R_Typ == 8'h1; // @[helpers.scala 65:24]
  assign _T_73 = output_[7]; // @[helpers.scala 65:51]
  assign _T_75 = _T_73 ? 24'hffffff : 24'h0; // @[Bitwise.scala 71:12]
  assign _T_76 = output_[7:0]; // @[helpers.scala 65:61]
  assign _T_77 = {_T_75,_T_76}; // @[Cat.scala 29:58]
  assign _T_78 = request_R_Typ == 8'h5; // @[helpers.scala 66:26]
  assign _T_81 = {24'h0,_T_76}; // @[Cat.scala 29:58]
  assign _T_83 = _T_78 ? _T_81 : output_; // @[helpers.scala 66:14]
  assign _T_84 = _T_72 ? _T_77 : _T_83; // @[helpers.scala 65:12]
  assign _T_85 = _T_68 ? _T_71 : _T_84; // @[helpers.scala 64:10]
  assign _T_86 = _T_62 ? _T_67 : _T_85; // @[helpers.scala 63:18]
  assign _GEN_21 = _T_56 ? _T_86 : 32'h0; // @[Conditional.scala 39:67]
  assign _GEN_30 = _T_52 ? 1'h0 : _T_56; // @[Conditional.scala 39:67]
  assign _GEN_32 = _T_52 ? 32'h0 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_50 ? _GEN_8 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_41 = _T_50 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_43 = _T_50 ? 32'h0 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_48 = _T_48 ? _GEN_6 : _GEN_36; // @[Conditional.scala 40:58]
  assign io_NodeReq_ready = state == 2'h0; // @[ReadMemoryController.scala 83:20]
  assign io_MemReq_valid = _T_48 ? 1'h0 : _T_50; // @[ReadMemoryController.scala 95:19 ReadMemoryController.scala 140:23]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_57; // @[ReadMemoryController.scala 96:23]
  assign io_MemReq_bits_tag = {{7'd0}, ID}; // @[ReadMemoryController.scala 99:22]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[ReadMemoryController.scala 104:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[ReadMemoryController.scala 101:26]
  assign io_output_valid = _T_48 ? 1'h0 : _GEN_41; // @[ReadMemoryController.scala 90:19 ReadMemoryController.scala 164:23]
  assign io_output_bits_RouteID = request_R_RouteID; // @[ReadMemoryController.scala 91:26]
  assign io_output_bits_data = _T_48 ? 32'h0 : _GEN_43; // @[ReadMemoryController.scala 93:23 ReadMemoryController.scala 168:29]
  assign io_free = state == 2'h0; // @[ReadMemoryController.scala 81:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ID = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_RouteID = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  request_R_address = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  request_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  request_R_Typ = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  bitmask = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sendbytemask = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ReqAddress = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ptr = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  linebuffer_0 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  linebuffer_1 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  isWrite = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    ID <= reset;
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_9) begin
        request_R_RouteID <= io_NodeReq_bits_RouteID;
      end
    end
    if (reset) begin
      request_R_address <= 32'h0;
    end else begin
      if (_T_9) begin
        request_R_address <= io_NodeReq_bits_address;
      end
    end
    if (reset) begin
      request_R_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      request_R_Typ <= 8'h3;
    end else begin
      if (_T_9) begin
        request_R_Typ <= io_NodeReq_bits_Typ;
      end
    end
    if (reset) begin
      bitmask <= 64'h0;
    end else begin
      bitmask <= _GEN_5[63:0];
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_48[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_9) begin
        ReqAddress <= _T_11;
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              ptr <= _T_54;
            end
          end else begin
            if (_T_56) begin
              ptr <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (1'h0 == ptr) begin
                linebuffer_0 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (ptr) begin
                linebuffer_1 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_48) begin
        if (_T_9) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_50) begin
          if (io_MemReq_ready) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (_T_55) begin
                state <= 2'h3;
              end else begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_56) begin
              if (io_output_ready) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    isWrite <= reset;
  end
endmodule
module ReadTableEntry_1(
  input         clock,
  input         reset,
  output        io_NodeReq_ready,
  input         io_NodeReq_valid,
  input  [15:0] io_NodeReq_bits_RouteID,
  input  [31:0] io_NodeReq_bits_address,
  input  [4:0]  io_NodeReq_bits_taskID,
  input  [7:0]  io_NodeReq_bits_Typ,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_data,
  input         io_output_ready,
  output        io_output_valid,
  output [15:0] io_output_bits_RouteID,
  output [31:0] io_output_bits_data,
  output        io_free
);
  reg  ID; // @[ReadMemoryController.scala 49:19]
  reg [31:0] _RAND_0;
  reg [15:0] request_R_RouteID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_1;
  reg [31:0] request_R_address; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_2;
  reg [4:0] request_R_taskID; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_3;
  reg [7:0] request_R_Typ; // @[ReadMemoryController.scala 51:32]
  reg [31:0] _RAND_4;
  reg [63:0] bitmask; // @[ReadMemoryController.scala 56:29]
  reg [63:0] _RAND_5;
  reg [7:0] sendbytemask; // @[ReadMemoryController.scala 58:29]
  reg [31:0] _RAND_6;
  reg [31:0] ReqAddress; // @[ReadMemoryController.scala 62:27]
  reg [31:0] _RAND_7;
  reg  ptr; // @[ReadMemoryController.scala 66:27]
  reg [31:0] _RAND_8;
  reg [31:0] linebuffer_0; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_9;
  reg [31:0] linebuffer_1; // @[ReadMemoryController.scala 67:27]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[ReadMemoryController.scala 73:68]
  reg [31:0] _RAND_11;
  wire [2:0] _T_6; // @[Cat.scala 29:58]
  wire [31:0] _GEN_57; // @[ReadMemoryController.scala 96:37]
  reg  isWrite; // @[ReadMemoryController.scala 100:24]
  reg [31:0] _RAND_12;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire [29:0] _T_10; // @[ReadMemoryController.scala 115:44]
  wire [31:0] _T_11; // @[ReadMemoryController.scala 115:69]
  wire  _T_12; // @[helpers.scala 27:24]
  wire  _T_13; // @[helpers.scala 27:47]
  wire  _T_14; // @[helpers.scala 27:40]
  wire  _T_16; // @[helpers.scala 28:15]
  wire  _T_17; // @[helpers.scala 28:38]
  wire  _T_18; // @[helpers.scala 28:31]
  wire  _T_20; // @[helpers.scala 29:17]
  wire  _T_21; // @[helpers.scala 29:40]
  wire  _T_22; // @[helpers.scala 29:33]
  wire [63:0] _T_25; // @[helpers.scala 29:12]
  wire [63:0] _T_26; // @[helpers.scala 28:10]
  wire [63:0] _T_27; // @[helpers.scala 27:19]
  wire [1:0] _T_28; // @[helpers.scala 39:32]
  wire [4:0] _T_29; // @[Cat.scala 29:58]
  wire [94:0] _GEN_58; // @[helpers.scala 40:26]
  wire [94:0] _T_30; // @[helpers.scala 40:26]
  wire [7:0] _T_43; // @[helpers.scala 50:12]
  wire [7:0] _T_44; // @[helpers.scala 49:10]
  wire [7:0] _T_45; // @[helpers.scala 48:19]
  wire [10:0] _GEN_59; // @[helpers.scala 20:26]
  wire [10:0] _T_47; // @[helpers.scala 20:26]
  wire [94:0] _GEN_5; // @[ReadMemoryController.scala 111:28]
  wire [10:0] _GEN_6; // @[ReadMemoryController.scala 111:28]
  wire  _T_48; // @[Conditional.scala 37:30]
  wire  _T_50; // @[Conditional.scala 37:30]
  wire [3:0] _T_51; // @[ReadMemoryController.scala 144:38]
  wire [10:0] _GEN_8; // @[ReadMemoryController.scala 142:29]
  wire  _T_52; // @[Conditional.scala 37:30]
  wire  _T_54; // @[ReadMemoryController.scala 154:20]
  wire  _T_55; // @[ReadMemoryController.scala 156:27]
  wire  _T_56; // @[Conditional.scala 37:30]
  wire [63:0] _T_57; // @[ReadMemoryController.scala 165:29]
  wire [63:0] _T_58; // @[ReadMemoryController.scala 165:36]
  wire [1:0] _T_59; // @[ReadMemoryController.scala 165:71]
  wire [4:0] _T_60; // @[Cat.scala 29:58]
  wire [63:0] _T_61; // @[ReadMemoryController.scala 165:47]
  wire  _T_62; // @[helpers.scala 63:30]
  wire [63:0] _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_31; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_42; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_53; // @[Conditional.scala 40:58]
  wire [31:0] output_; // @[ReadMemoryController.scala 165:14]
  wire  _T_63; // @[helpers.scala 63:57]
  wire [15:0] _T_65; // @[Bitwise.scala 71:12]
  wire [15:0] _T_66; // @[helpers.scala 63:68]
  wire [31:0] _T_67; // @[Cat.scala 29:58]
  wire  _T_68; // @[helpers.scala 64:22]
  wire [31:0] _T_71; // @[Cat.scala 29:58]
  wire  _T_72; // @[helpers.scala 65:24]
  wire  _T_73; // @[helpers.scala 65:51]
  wire [23:0] _T_75; // @[Bitwise.scala 71:12]
  wire [7:0] _T_76; // @[helpers.scala 65:61]
  wire [31:0] _T_77; // @[Cat.scala 29:58]
  wire  _T_78; // @[helpers.scala 66:26]
  wire [31:0] _T_81; // @[Cat.scala 29:58]
  wire [31:0] _T_83; // @[helpers.scala 66:14]
  wire [31:0] _T_84; // @[helpers.scala 65:12]
  wire [31:0] _T_85; // @[helpers.scala 64:10]
  wire [31:0] _T_86; // @[helpers.scala 63:18]
  wire [31:0] _GEN_21; // @[Conditional.scala 39:67]
  wire  _GEN_30; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_32; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_41; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_43; // @[Conditional.scala 39:67]
  wire [10:0] _GEN_48; // @[Conditional.scala 40:58]
  assign _T_6 = {ptr,2'h0}; // @[Cat.scala 29:58]
  assign _GEN_57 = {{29'd0}, _T_6}; // @[ReadMemoryController.scala 96:37]
  assign _T_9 = io_NodeReq_ready & io_NodeReq_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_NodeReq_bits_address[31:2]; // @[ReadMemoryController.scala 115:44]
  assign _T_11 = {_T_10, 2'h0}; // @[ReadMemoryController.scala 115:69]
  assign _T_12 = io_NodeReq_bits_Typ == 8'h2; // @[helpers.scala 27:24]
  assign _T_13 = io_NodeReq_bits_Typ == 8'h6; // @[helpers.scala 27:47]
  assign _T_14 = _T_12 | _T_13; // @[helpers.scala 27:40]
  assign _T_16 = io_NodeReq_bits_Typ == 8'h1; // @[helpers.scala 28:15]
  assign _T_17 = io_NodeReq_bits_Typ == 8'h5; // @[helpers.scala 28:38]
  assign _T_18 = _T_16 | _T_17; // @[helpers.scala 28:31]
  assign _T_20 = io_NodeReq_bits_Typ == 8'h3; // @[helpers.scala 29:17]
  assign _T_21 = io_NodeReq_bits_Typ == 8'h7; // @[helpers.scala 29:40]
  assign _T_22 = _T_20 | _T_21; // @[helpers.scala 29:33]
  assign _T_25 = _T_22 ? 64'hffffffff : 64'hffffffffffffffff; // @[helpers.scala 29:12]
  assign _T_26 = _T_18 ? 64'hff : _T_25; // @[helpers.scala 28:10]
  assign _T_27 = _T_14 ? 64'hffff : _T_26; // @[helpers.scala 27:19]
  assign _T_28 = io_NodeReq_bits_address[1:0]; // @[helpers.scala 39:32]
  assign _T_29 = {_T_28,3'h0}; // @[Cat.scala 29:58]
  assign _GEN_58 = {{31'd0}, _T_27}; // @[helpers.scala 40:26]
  assign _T_30 = _GEN_58 << _T_29; // @[helpers.scala 40:26]
  assign _T_43 = _T_22 ? 8'hf : 8'hff; // @[helpers.scala 50:12]
  assign _T_44 = _T_18 ? 8'h1 : _T_43; // @[helpers.scala 49:10]
  assign _T_45 = _T_14 ? 8'h3 : _T_44; // @[helpers.scala 48:19]
  assign _GEN_59 = {{3'd0}, _T_45}; // @[helpers.scala 20:26]
  assign _T_47 = _GEN_59 << _T_28; // @[helpers.scala 20:26]
  assign _GEN_5 = _T_9 ? _T_30 : {{31'd0}, bitmask}; // @[ReadMemoryController.scala 111:28]
  assign _GEN_6 = _T_9 ? _T_47 : {{3'd0}, sendbytemask}; // @[ReadMemoryController.scala 111:28]
  assign _T_48 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_50 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_51 = sendbytemask[7:4]; // @[ReadMemoryController.scala 144:38]
  assign _GEN_8 = io_MemReq_ready ? {{7'd0}, _T_51} : _GEN_6; // @[ReadMemoryController.scala 142:29]
  assign _T_52 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_54 = ptr + 1'h1; // @[ReadMemoryController.scala 154:20]
  assign _T_55 = sendbytemask == 8'h0; // @[ReadMemoryController.scala 156:27]
  assign _T_56 = 2'h3 == state; // @[Conditional.scala 37:30]
  assign _T_57 = {linebuffer_1,linebuffer_0}; // @[ReadMemoryController.scala 165:29]
  assign _T_58 = _T_57 & bitmask; // @[ReadMemoryController.scala 165:36]
  assign _T_59 = request_R_address[1:0]; // @[ReadMemoryController.scala 165:71]
  assign _T_60 = {_T_59,3'h0}; // @[Cat.scala 29:58]
  assign _T_61 = _T_58 >> _T_60; // @[ReadMemoryController.scala 165:47]
  assign _T_62 = request_R_Typ == 8'h2; // @[helpers.scala 63:30]
  assign _GEN_20 = _T_56 ? _T_61 : 64'h0; // @[Conditional.scala 39:67]
  assign _GEN_31 = _T_52 ? 64'h0 : _GEN_20; // @[Conditional.scala 39:67]
  assign _GEN_42 = _T_50 ? 64'h0 : _GEN_31; // @[Conditional.scala 39:67]
  assign _GEN_53 = _T_48 ? 64'h0 : _GEN_42; // @[Conditional.scala 40:58]
  assign output_ = _GEN_53[31:0]; // @[ReadMemoryController.scala 165:14]
  assign _T_63 = output_[15]; // @[helpers.scala 63:57]
  assign _T_65 = _T_63 ? 16'hffff : 16'h0; // @[Bitwise.scala 71:12]
  assign _T_66 = output_[15:0]; // @[helpers.scala 63:68]
  assign _T_67 = {_T_65,_T_66}; // @[Cat.scala 29:58]
  assign _T_68 = request_R_Typ == 8'h6; // @[helpers.scala 64:22]
  assign _T_71 = {16'h0,_T_66}; // @[Cat.scala 29:58]
  assign _T_72 = request_R_Typ == 8'h1; // @[helpers.scala 65:24]
  assign _T_73 = output_[7]; // @[helpers.scala 65:51]
  assign _T_75 = _T_73 ? 24'hffffff : 24'h0; // @[Bitwise.scala 71:12]
  assign _T_76 = output_[7:0]; // @[helpers.scala 65:61]
  assign _T_77 = {_T_75,_T_76}; // @[Cat.scala 29:58]
  assign _T_78 = request_R_Typ == 8'h5; // @[helpers.scala 66:26]
  assign _T_81 = {24'h0,_T_76}; // @[Cat.scala 29:58]
  assign _T_83 = _T_78 ? _T_81 : output_; // @[helpers.scala 66:14]
  assign _T_84 = _T_72 ? _T_77 : _T_83; // @[helpers.scala 65:12]
  assign _T_85 = _T_68 ? _T_71 : _T_84; // @[helpers.scala 64:10]
  assign _T_86 = _T_62 ? _T_67 : _T_85; // @[helpers.scala 63:18]
  assign _GEN_21 = _T_56 ? _T_86 : 32'h0; // @[Conditional.scala 39:67]
  assign _GEN_30 = _T_52 ? 1'h0 : _T_56; // @[Conditional.scala 39:67]
  assign _GEN_32 = _T_52 ? 32'h0 : _GEN_21; // @[Conditional.scala 39:67]
  assign _GEN_36 = _T_50 ? _GEN_8 : _GEN_6; // @[Conditional.scala 39:67]
  assign _GEN_41 = _T_50 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67]
  assign _GEN_43 = _T_50 ? 32'h0 : _GEN_32; // @[Conditional.scala 39:67]
  assign _GEN_48 = _T_48 ? _GEN_6 : _GEN_36; // @[Conditional.scala 40:58]
  assign io_NodeReq_ready = state == 2'h0; // @[ReadMemoryController.scala 83:20]
  assign io_MemReq_valid = _T_48 ? 1'h0 : _T_50; // @[ReadMemoryController.scala 95:19 ReadMemoryController.scala 140:23]
  assign io_MemReq_bits_addr = ReqAddress + _GEN_57; // @[ReadMemoryController.scala 96:23]
  assign io_MemReq_bits_tag = {{7'd0}, ID}; // @[ReadMemoryController.scala 99:22]
  assign io_MemReq_bits_taskID = request_R_taskID; // @[ReadMemoryController.scala 104:25]
  assign io_MemReq_bits_iswrite = isWrite; // @[ReadMemoryController.scala 101:26]
  assign io_output_valid = _T_48 ? 1'h0 : _GEN_41; // @[ReadMemoryController.scala 90:19 ReadMemoryController.scala 164:23]
  assign io_output_bits_RouteID = request_R_RouteID; // @[ReadMemoryController.scala 91:26]
  assign io_output_bits_data = _T_48 ? 32'h0 : _GEN_43; // @[ReadMemoryController.scala 93:23 ReadMemoryController.scala 168:29]
  assign io_free = state == 2'h0; // @[ReadMemoryController.scala 81:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ID = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  request_R_RouteID = _RAND_1[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  request_R_address = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  request_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  request_R_Typ = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  bitmask = _RAND_5[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  sendbytemask = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ReqAddress = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ptr = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  linebuffer_0 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  linebuffer_1 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  isWrite = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      ID <= 1'h0;
    end else begin
      ID <= 1'h1;
    end
    if (reset) begin
      request_R_RouteID <= 16'h0;
    end else begin
      if (_T_9) begin
        request_R_RouteID <= io_NodeReq_bits_RouteID;
      end
    end
    if (reset) begin
      request_R_address <= 32'h0;
    end else begin
      if (_T_9) begin
        request_R_address <= io_NodeReq_bits_address;
      end
    end
    if (reset) begin
      request_R_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        request_R_taskID <= io_NodeReq_bits_taskID;
      end
    end
    if (reset) begin
      request_R_Typ <= 8'h3;
    end else begin
      if (_T_9) begin
        request_R_Typ <= io_NodeReq_bits_Typ;
      end
    end
    if (reset) begin
      bitmask <= 64'h0;
    end else begin
      bitmask <= _GEN_5[63:0];
    end
    if (reset) begin
      sendbytemask <= 8'h0;
    end else begin
      sendbytemask <= _GEN_48[7:0];
    end
    if (reset) begin
      ReqAddress <= 32'h0;
    end else begin
      if (_T_9) begin
        ReqAddress <= _T_11;
      end
    end
    if (reset) begin
      ptr <= 1'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              ptr <= _T_54;
            end
          end else begin
            if (_T_56) begin
              ptr <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_0 <= 32'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (1'h0 == ptr) begin
                linebuffer_0 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      linebuffer_1 <= 32'h0;
    end else begin
      if (!(_T_48)) begin
        if (!(_T_50)) begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (ptr) begin
                linebuffer_1 <= io_MemResp_data;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_48) begin
        if (_T_9) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_50) begin
          if (io_MemReq_ready) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_52) begin
            if (io_MemResp_valid) begin
              if (_T_55) begin
                state <= 2'h3;
              end else begin
                state <= 2'h1;
              end
            end
          end else begin
            if (_T_56) begin
              if (io_output_ready) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    isWrite <= reset;
  end
endmodule
module ReadMemoryController(
  input         clock,
  input         reset,
  output        io_ReadIn_0_ready,
  input         io_ReadIn_0_valid,
  input  [31:0] io_ReadIn_0_bits_address,
  input  [4:0]  io_ReadIn_0_bits_taskID,
  output        io_ReadIn_1_ready,
  input         io_ReadIn_1_valid,
  input  [31:0] io_ReadIn_1_bits_address,
  input  [4:0]  io_ReadIn_1_bits_taskID,
  output        io_ReadIn_2_ready,
  input         io_ReadIn_2_valid,
  input  [31:0] io_ReadIn_2_bits_address,
  input  [4:0]  io_ReadIn_2_bits_taskID,
  output        io_ReadIn_3_ready,
  input         io_ReadIn_3_valid,
  input  [31:0] io_ReadIn_3_bits_address,
  input  [4:0]  io_ReadIn_3_bits_taskID,
  output        io_ReadIn_4_ready,
  input         io_ReadIn_4_valid,
  input  [31:0] io_ReadIn_4_bits_address,
  input  [4:0]  io_ReadIn_4_bits_taskID,
  output        io_ReadIn_5_ready,
  input         io_ReadIn_5_valid,
  input  [31:0] io_ReadIn_5_bits_address,
  input  [4:0]  io_ReadIn_5_bits_taskID,
  output        io_ReadIn_6_ready,
  input         io_ReadIn_6_valid,
  input  [31:0] io_ReadIn_6_bits_address,
  input  [4:0]  io_ReadIn_6_bits_taskID,
  output        io_ReadIn_7_ready,
  input         io_ReadIn_7_valid,
  input  [31:0] io_ReadIn_7_bits_address,
  input  [4:0]  io_ReadIn_7_bits_taskID,
  output        io_ReadIn_8_ready,
  input         io_ReadIn_8_valid,
  input  [31:0] io_ReadIn_8_bits_address,
  input  [4:0]  io_ReadIn_8_bits_taskID,
  output        io_ReadIn_9_ready,
  input         io_ReadIn_9_valid,
  input  [31:0] io_ReadIn_9_bits_address,
  input  [4:0]  io_ReadIn_9_bits_taskID,
  output        io_ReadIn_10_ready,
  input         io_ReadIn_10_valid,
  input  [31:0] io_ReadIn_10_bits_address,
  input  [4:0]  io_ReadIn_10_bits_taskID,
  output        io_ReadIn_11_ready,
  input         io_ReadIn_11_valid,
  input  [31:0] io_ReadIn_11_bits_address,
  input  [4:0]  io_ReadIn_11_bits_taskID,
  output        io_ReadIn_12_ready,
  input         io_ReadIn_12_valid,
  input  [31:0] io_ReadIn_12_bits_address,
  input  [4:0]  io_ReadIn_12_bits_taskID,
  output        io_ReadIn_13_ready,
  input         io_ReadIn_13_valid,
  input  [31:0] io_ReadIn_13_bits_address,
  input  [4:0]  io_ReadIn_13_bits_taskID,
  output        io_ReadIn_14_ready,
  input         io_ReadIn_14_valid,
  input  [31:0] io_ReadIn_14_bits_address,
  input  [4:0]  io_ReadIn_14_bits_taskID,
  output        io_ReadIn_15_ready,
  input         io_ReadIn_15_valid,
  input  [31:0] io_ReadIn_15_bits_address,
  input  [4:0]  io_ReadIn_15_bits_taskID,
  output        io_ReadIn_16_ready,
  input         io_ReadIn_16_valid,
  input  [31:0] io_ReadIn_16_bits_address,
  input  [4:0]  io_ReadIn_16_bits_taskID,
  output        io_ReadIn_17_ready,
  input         io_ReadIn_17_valid,
  input  [31:0] io_ReadIn_17_bits_address,
  input  [4:0]  io_ReadIn_17_bits_taskID,
  output        io_ReadIn_18_ready,
  input         io_ReadIn_18_valid,
  input  [31:0] io_ReadIn_18_bits_address,
  input  [4:0]  io_ReadIn_18_bits_taskID,
  output        io_ReadOut_0_valid,
  output [31:0] io_ReadOut_0_data,
  output        io_ReadOut_1_valid,
  output [31:0] io_ReadOut_1_data,
  output        io_ReadOut_2_valid,
  output [31:0] io_ReadOut_2_data,
  output        io_ReadOut_3_valid,
  output [31:0] io_ReadOut_3_data,
  output        io_ReadOut_4_valid,
  output [31:0] io_ReadOut_4_data,
  output        io_ReadOut_5_valid,
  output [31:0] io_ReadOut_5_data,
  output        io_ReadOut_6_valid,
  output [31:0] io_ReadOut_6_data,
  output        io_ReadOut_7_valid,
  output [31:0] io_ReadOut_7_data,
  output        io_ReadOut_8_valid,
  output [31:0] io_ReadOut_8_data,
  output        io_ReadOut_9_valid,
  output [31:0] io_ReadOut_9_data,
  output        io_ReadOut_10_valid,
  output [31:0] io_ReadOut_10_data,
  output        io_ReadOut_11_valid,
  output [31:0] io_ReadOut_11_data,
  output        io_ReadOut_12_valid,
  output [31:0] io_ReadOut_12_data,
  output        io_ReadOut_13_valid,
  output [31:0] io_ReadOut_13_data,
  output        io_ReadOut_14_valid,
  output [31:0] io_ReadOut_14_data,
  output        io_ReadOut_15_valid,
  output [31:0] io_ReadOut_15_data,
  output        io_ReadOut_16_valid,
  output [31:0] io_ReadOut_16_data,
  output        io_ReadOut_17_valid,
  output [31:0] io_ReadOut_17_data,
  output        io_ReadOut_18_valid,
  output [31:0] io_ReadOut_18_data,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag
);
  wire  in_arb_clock; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_0_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_0_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_0_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_0_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_1_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_1_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_1_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_1_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_2_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_2_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_2_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_2_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_3_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_3_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_3_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_3_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_4_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_4_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_4_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_4_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_5_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_5_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_5_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_5_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_6_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_6_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_6_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_6_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_7_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_7_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_7_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_7_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_8_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_8_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_8_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_8_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_9_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_9_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_9_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_9_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_10_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_10_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_10_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_10_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_11_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_11_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_11_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_11_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_12_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_12_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_12_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_12_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_13_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_13_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_13_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_13_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_14_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_14_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_14_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_14_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_15_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_15_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_15_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_15_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_16_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_16_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_16_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_16_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_17_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_17_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_17_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_17_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_18_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_in_18_valid; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_in_18_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_in_18_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_out_ready; // @[ReadMemoryController.scala 221:25]
  wire  in_arb_io_out_valid; // @[ReadMemoryController.scala 221:25]
  wire [15:0] in_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 221:25]
  wire [31:0] in_arb_io_out_bits_address; // @[ReadMemoryController.scala 221:25]
  wire [4:0] in_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 221:25]
  wire [7:0] in_arb_io_out_bits_Typ; // @[ReadMemoryController.scala 221:25]
  wire  alloc_arb_io_in_0_ready; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_in_0_valid; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_in_1_ready; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_in_1_valid; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_out_ready; // @[ReadMemoryController.scala 223:25]
  wire  alloc_arb_io_out_valid; // @[ReadMemoryController.scala 223:25]
  wire  cachereq_arb_io_in_0_ready; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_0_valid; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_0_bits_addr; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_0_bits_data; // @[ReadMemoryController.scala 226:31]
  wire [3:0] cachereq_arb_io_in_0_bits_mask; // @[ReadMemoryController.scala 226:31]
  wire [7:0] cachereq_arb_io_in_0_bits_tag; // @[ReadMemoryController.scala 226:31]
  wire [4:0] cachereq_arb_io_in_0_bits_taskID; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_0_bits_iswrite; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_1_ready; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_1_valid; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_1_bits_addr; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_in_1_bits_data; // @[ReadMemoryController.scala 226:31]
  wire [3:0] cachereq_arb_io_in_1_bits_mask; // @[ReadMemoryController.scala 226:31]
  wire [7:0] cachereq_arb_io_in_1_bits_tag; // @[ReadMemoryController.scala 226:31]
  wire [4:0] cachereq_arb_io_in_1_bits_taskID; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_in_1_bits_iswrite; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_out_ready; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_out_valid; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_out_bits_addr; // @[ReadMemoryController.scala 226:31]
  wire [31:0] cachereq_arb_io_out_bits_data; // @[ReadMemoryController.scala 226:31]
  wire [3:0] cachereq_arb_io_out_bits_mask; // @[ReadMemoryController.scala 226:31]
  wire [7:0] cachereq_arb_io_out_bits_tag; // @[ReadMemoryController.scala 226:31]
  wire [4:0] cachereq_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 226:31]
  wire  cachereq_arb_io_out_bits_iswrite; // @[ReadMemoryController.scala 226:31]
  wire  cacheresp_demux_io_en; // @[ReadMemoryController.scala 228:31]
  wire [31:0] cacheresp_demux_io_input_data; // @[ReadMemoryController.scala 228:31]
  wire [7:0] cacheresp_demux_io_input_tag; // @[ReadMemoryController.scala 228:31]
  wire  cacheresp_demux_io_sel; // @[ReadMemoryController.scala 228:31]
  wire  cacheresp_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 228:31]
  wire [31:0] cacheresp_demux_io_outputs_0_data; // @[ReadMemoryController.scala 228:31]
  wire [7:0] cacheresp_demux_io_outputs_0_tag; // @[ReadMemoryController.scala 228:31]
  wire  cacheresp_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 228:31]
  wire [31:0] cacheresp_demux_io_outputs_1_data; // @[ReadMemoryController.scala 228:31]
  wire [7:0] cacheresp_demux_io_outputs_1_tag; // @[ReadMemoryController.scala 228:31]
  wire  out_arb_clock; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_0_ready; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_0_valid; // @[ReadMemoryController.scala 231:25]
  wire [15:0] out_arb_io_in_0_bits_RouteID; // @[ReadMemoryController.scala 231:25]
  wire [31:0] out_arb_io_in_0_bits_data; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_1_ready; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_in_1_valid; // @[ReadMemoryController.scala 231:25]
  wire [15:0] out_arb_io_in_1_bits_RouteID; // @[ReadMemoryController.scala 231:25]
  wire [31:0] out_arb_io_in_1_bits_data; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_out_ready; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_out_valid; // @[ReadMemoryController.scala 231:25]
  wire [15:0] out_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 231:25]
  wire [31:0] out_arb_io_out_bits_data; // @[ReadMemoryController.scala 231:25]
  wire  out_arb_io_chosen; // @[ReadMemoryController.scala 231:25]
  wire  out_demux_clock; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_reset; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_0_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_1_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_2_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_2_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_3_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_3_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_4_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_4_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_5_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_5_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_6_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_6_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_7_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_7_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_8_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_8_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_9_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_9_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_10_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_10_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_11_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_11_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_12_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_12_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_13_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_13_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_14_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_14_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_15_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_15_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_16_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_16_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_17_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_17_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_outputs_18_valid; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_outputs_18_data; // @[ReadMemoryController.scala 232:25]
  wire [15:0] out_demux_io_input_RouteID; // @[ReadMemoryController.scala 232:25]
  wire [31:0] out_demux_io_input_data; // @[ReadMemoryController.scala 232:25]
  wire  out_demux_io_enable; // @[ReadMemoryController.scala 232:25]
  wire  ReadTable_0_clock; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_reset; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_NodeReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_NodeReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_0_io_NodeReq_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_NodeReq_bits_address; // @[ReadMemoryController.scala 251:28]
  wire [4:0] ReadTable_0_io_NodeReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_0_io_NodeReq_bits_Typ; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_MemReq_bits_addr; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_0_io_MemReq_bits_tag; // @[ReadMemoryController.scala 251:28]
  wire [4:0] ReadTable_0_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_MemResp_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_MemResp_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_output_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_output_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_0_io_output_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_0_io_output_bits_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_0_io_free; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_clock; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_reset; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_NodeReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_NodeReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_1_io_NodeReq_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_NodeReq_bits_address; // @[ReadMemoryController.scala 251:28]
  wire [4:0] ReadTable_1_io_NodeReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_1_io_NodeReq_bits_Typ; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemReq_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemReq_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_MemReq_bits_addr; // @[ReadMemoryController.scala 251:28]
  wire [7:0] ReadTable_1_io_MemReq_bits_tag; // @[ReadMemoryController.scala 251:28]
  wire [4:0] ReadTable_1_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_MemResp_valid; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_MemResp_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_output_ready; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_output_valid; // @[ReadMemoryController.scala 251:28]
  wire [15:0] ReadTable_1_io_output_bits_RouteID; // @[ReadMemoryController.scala 251:28]
  wire [31:0] ReadTable_1_io_output_bits_data; // @[ReadMemoryController.scala 251:28]
  wire  ReadTable_1_io_free; // @[ReadMemoryController.scala 251:28]
  ArbiterTree_1 in_arb ( // @[ReadMemoryController.scala 221:25]
    .clock(in_arb_clock),
    .io_in_0_ready(in_arb_io_in_0_ready),
    .io_in_0_valid(in_arb_io_in_0_valid),
    .io_in_0_bits_address(in_arb_io_in_0_bits_address),
    .io_in_0_bits_taskID(in_arb_io_in_0_bits_taskID),
    .io_in_1_ready(in_arb_io_in_1_ready),
    .io_in_1_valid(in_arb_io_in_1_valid),
    .io_in_1_bits_address(in_arb_io_in_1_bits_address),
    .io_in_1_bits_taskID(in_arb_io_in_1_bits_taskID),
    .io_in_2_ready(in_arb_io_in_2_ready),
    .io_in_2_valid(in_arb_io_in_2_valid),
    .io_in_2_bits_address(in_arb_io_in_2_bits_address),
    .io_in_2_bits_taskID(in_arb_io_in_2_bits_taskID),
    .io_in_3_ready(in_arb_io_in_3_ready),
    .io_in_3_valid(in_arb_io_in_3_valid),
    .io_in_3_bits_address(in_arb_io_in_3_bits_address),
    .io_in_3_bits_taskID(in_arb_io_in_3_bits_taskID),
    .io_in_4_ready(in_arb_io_in_4_ready),
    .io_in_4_valid(in_arb_io_in_4_valid),
    .io_in_4_bits_address(in_arb_io_in_4_bits_address),
    .io_in_4_bits_taskID(in_arb_io_in_4_bits_taskID),
    .io_in_5_ready(in_arb_io_in_5_ready),
    .io_in_5_valid(in_arb_io_in_5_valid),
    .io_in_5_bits_address(in_arb_io_in_5_bits_address),
    .io_in_5_bits_taskID(in_arb_io_in_5_bits_taskID),
    .io_in_6_ready(in_arb_io_in_6_ready),
    .io_in_6_valid(in_arb_io_in_6_valid),
    .io_in_6_bits_address(in_arb_io_in_6_bits_address),
    .io_in_6_bits_taskID(in_arb_io_in_6_bits_taskID),
    .io_in_7_ready(in_arb_io_in_7_ready),
    .io_in_7_valid(in_arb_io_in_7_valid),
    .io_in_7_bits_address(in_arb_io_in_7_bits_address),
    .io_in_7_bits_taskID(in_arb_io_in_7_bits_taskID),
    .io_in_8_ready(in_arb_io_in_8_ready),
    .io_in_8_valid(in_arb_io_in_8_valid),
    .io_in_8_bits_address(in_arb_io_in_8_bits_address),
    .io_in_8_bits_taskID(in_arb_io_in_8_bits_taskID),
    .io_in_9_ready(in_arb_io_in_9_ready),
    .io_in_9_valid(in_arb_io_in_9_valid),
    .io_in_9_bits_address(in_arb_io_in_9_bits_address),
    .io_in_9_bits_taskID(in_arb_io_in_9_bits_taskID),
    .io_in_10_ready(in_arb_io_in_10_ready),
    .io_in_10_valid(in_arb_io_in_10_valid),
    .io_in_10_bits_address(in_arb_io_in_10_bits_address),
    .io_in_10_bits_taskID(in_arb_io_in_10_bits_taskID),
    .io_in_11_ready(in_arb_io_in_11_ready),
    .io_in_11_valid(in_arb_io_in_11_valid),
    .io_in_11_bits_address(in_arb_io_in_11_bits_address),
    .io_in_11_bits_taskID(in_arb_io_in_11_bits_taskID),
    .io_in_12_ready(in_arb_io_in_12_ready),
    .io_in_12_valid(in_arb_io_in_12_valid),
    .io_in_12_bits_address(in_arb_io_in_12_bits_address),
    .io_in_12_bits_taskID(in_arb_io_in_12_bits_taskID),
    .io_in_13_ready(in_arb_io_in_13_ready),
    .io_in_13_valid(in_arb_io_in_13_valid),
    .io_in_13_bits_address(in_arb_io_in_13_bits_address),
    .io_in_13_bits_taskID(in_arb_io_in_13_bits_taskID),
    .io_in_14_ready(in_arb_io_in_14_ready),
    .io_in_14_valid(in_arb_io_in_14_valid),
    .io_in_14_bits_address(in_arb_io_in_14_bits_address),
    .io_in_14_bits_taskID(in_arb_io_in_14_bits_taskID),
    .io_in_15_ready(in_arb_io_in_15_ready),
    .io_in_15_valid(in_arb_io_in_15_valid),
    .io_in_15_bits_address(in_arb_io_in_15_bits_address),
    .io_in_15_bits_taskID(in_arb_io_in_15_bits_taskID),
    .io_in_16_ready(in_arb_io_in_16_ready),
    .io_in_16_valid(in_arb_io_in_16_valid),
    .io_in_16_bits_address(in_arb_io_in_16_bits_address),
    .io_in_16_bits_taskID(in_arb_io_in_16_bits_taskID),
    .io_in_17_ready(in_arb_io_in_17_ready),
    .io_in_17_valid(in_arb_io_in_17_valid),
    .io_in_17_bits_address(in_arb_io_in_17_bits_address),
    .io_in_17_bits_taskID(in_arb_io_in_17_bits_taskID),
    .io_in_18_ready(in_arb_io_in_18_ready),
    .io_in_18_valid(in_arb_io_in_18_valid),
    .io_in_18_bits_address(in_arb_io_in_18_bits_address),
    .io_in_18_bits_taskID(in_arb_io_in_18_bits_taskID),
    .io_out_ready(in_arb_io_out_ready),
    .io_out_valid(in_arb_io_out_valid),
    .io_out_bits_RouteID(in_arb_io_out_bits_RouteID),
    .io_out_bits_address(in_arb_io_out_bits_address),
    .io_out_bits_taskID(in_arb_io_out_bits_taskID),
    .io_out_bits_Typ(in_arb_io_out_bits_Typ)
  );
  Arbiter alloc_arb ( // @[ReadMemoryController.scala 223:25]
    .io_in_0_ready(alloc_arb_io_in_0_ready),
    .io_in_0_valid(alloc_arb_io_in_0_valid),
    .io_in_1_ready(alloc_arb_io_in_1_ready),
    .io_in_1_valid(alloc_arb_io_in_1_valid),
    .io_out_ready(alloc_arb_io_out_ready),
    .io_out_valid(alloc_arb_io_out_valid)
  );
  Arbiter_1 cachereq_arb ( // @[ReadMemoryController.scala 226:31]
    .io_in_0_ready(cachereq_arb_io_in_0_ready),
    .io_in_0_valid(cachereq_arb_io_in_0_valid),
    .io_in_0_bits_addr(cachereq_arb_io_in_0_bits_addr),
    .io_in_0_bits_data(cachereq_arb_io_in_0_bits_data),
    .io_in_0_bits_mask(cachereq_arb_io_in_0_bits_mask),
    .io_in_0_bits_tag(cachereq_arb_io_in_0_bits_tag),
    .io_in_0_bits_taskID(cachereq_arb_io_in_0_bits_taskID),
    .io_in_0_bits_iswrite(cachereq_arb_io_in_0_bits_iswrite),
    .io_in_1_ready(cachereq_arb_io_in_1_ready),
    .io_in_1_valid(cachereq_arb_io_in_1_valid),
    .io_in_1_bits_addr(cachereq_arb_io_in_1_bits_addr),
    .io_in_1_bits_data(cachereq_arb_io_in_1_bits_data),
    .io_in_1_bits_mask(cachereq_arb_io_in_1_bits_mask),
    .io_in_1_bits_tag(cachereq_arb_io_in_1_bits_tag),
    .io_in_1_bits_taskID(cachereq_arb_io_in_1_bits_taskID),
    .io_in_1_bits_iswrite(cachereq_arb_io_in_1_bits_iswrite),
    .io_out_ready(cachereq_arb_io_out_ready),
    .io_out_valid(cachereq_arb_io_out_valid),
    .io_out_bits_addr(cachereq_arb_io_out_bits_addr),
    .io_out_bits_data(cachereq_arb_io_out_bits_data),
    .io_out_bits_mask(cachereq_arb_io_out_bits_mask),
    .io_out_bits_tag(cachereq_arb_io_out_bits_tag),
    .io_out_bits_taskID(cachereq_arb_io_out_bits_taskID),
    .io_out_bits_iswrite(cachereq_arb_io_out_bits_iswrite)
  );
  Demux cacheresp_demux ( // @[ReadMemoryController.scala 228:31]
    .io_en(cacheresp_demux_io_en),
    .io_input_data(cacheresp_demux_io_input_data),
    .io_input_tag(cacheresp_demux_io_input_tag),
    .io_sel(cacheresp_demux_io_sel),
    .io_outputs_0_valid(cacheresp_demux_io_outputs_0_valid),
    .io_outputs_0_data(cacheresp_demux_io_outputs_0_data),
    .io_outputs_0_tag(cacheresp_demux_io_outputs_0_tag),
    .io_outputs_1_valid(cacheresp_demux_io_outputs_1_valid),
    .io_outputs_1_data(cacheresp_demux_io_outputs_1_data),
    .io_outputs_1_tag(cacheresp_demux_io_outputs_1_tag)
  );
  RRArbiter_1 out_arb ( // @[ReadMemoryController.scala 231:25]
    .clock(out_arb_clock),
    .io_in_0_ready(out_arb_io_in_0_ready),
    .io_in_0_valid(out_arb_io_in_0_valid),
    .io_in_0_bits_RouteID(out_arb_io_in_0_bits_RouteID),
    .io_in_0_bits_data(out_arb_io_in_0_bits_data),
    .io_in_1_ready(out_arb_io_in_1_ready),
    .io_in_1_valid(out_arb_io_in_1_valid),
    .io_in_1_bits_RouteID(out_arb_io_in_1_bits_RouteID),
    .io_in_1_bits_data(out_arb_io_in_1_bits_data),
    .io_out_ready(out_arb_io_out_ready),
    .io_out_valid(out_arb_io_out_valid),
    .io_out_bits_RouteID(out_arb_io_out_bits_RouteID),
    .io_out_bits_data(out_arb_io_out_bits_data),
    .io_chosen(out_arb_io_chosen)
  );
  DeMuxTree_1 out_demux ( // @[ReadMemoryController.scala 232:25]
    .clock(out_demux_clock),
    .reset(out_demux_reset),
    .io_outputs_0_valid(out_demux_io_outputs_0_valid),
    .io_outputs_0_data(out_demux_io_outputs_0_data),
    .io_outputs_1_valid(out_demux_io_outputs_1_valid),
    .io_outputs_1_data(out_demux_io_outputs_1_data),
    .io_outputs_2_valid(out_demux_io_outputs_2_valid),
    .io_outputs_2_data(out_demux_io_outputs_2_data),
    .io_outputs_3_valid(out_demux_io_outputs_3_valid),
    .io_outputs_3_data(out_demux_io_outputs_3_data),
    .io_outputs_4_valid(out_demux_io_outputs_4_valid),
    .io_outputs_4_data(out_demux_io_outputs_4_data),
    .io_outputs_5_valid(out_demux_io_outputs_5_valid),
    .io_outputs_5_data(out_demux_io_outputs_5_data),
    .io_outputs_6_valid(out_demux_io_outputs_6_valid),
    .io_outputs_6_data(out_demux_io_outputs_6_data),
    .io_outputs_7_valid(out_demux_io_outputs_7_valid),
    .io_outputs_7_data(out_demux_io_outputs_7_data),
    .io_outputs_8_valid(out_demux_io_outputs_8_valid),
    .io_outputs_8_data(out_demux_io_outputs_8_data),
    .io_outputs_9_valid(out_demux_io_outputs_9_valid),
    .io_outputs_9_data(out_demux_io_outputs_9_data),
    .io_outputs_10_valid(out_demux_io_outputs_10_valid),
    .io_outputs_10_data(out_demux_io_outputs_10_data),
    .io_outputs_11_valid(out_demux_io_outputs_11_valid),
    .io_outputs_11_data(out_demux_io_outputs_11_data),
    .io_outputs_12_valid(out_demux_io_outputs_12_valid),
    .io_outputs_12_data(out_demux_io_outputs_12_data),
    .io_outputs_13_valid(out_demux_io_outputs_13_valid),
    .io_outputs_13_data(out_demux_io_outputs_13_data),
    .io_outputs_14_valid(out_demux_io_outputs_14_valid),
    .io_outputs_14_data(out_demux_io_outputs_14_data),
    .io_outputs_15_valid(out_demux_io_outputs_15_valid),
    .io_outputs_15_data(out_demux_io_outputs_15_data),
    .io_outputs_16_valid(out_demux_io_outputs_16_valid),
    .io_outputs_16_data(out_demux_io_outputs_16_data),
    .io_outputs_17_valid(out_demux_io_outputs_17_valid),
    .io_outputs_17_data(out_demux_io_outputs_17_data),
    .io_outputs_18_valid(out_demux_io_outputs_18_valid),
    .io_outputs_18_data(out_demux_io_outputs_18_data),
    .io_input_RouteID(out_demux_io_input_RouteID),
    .io_input_data(out_demux_io_input_data),
    .io_enable(out_demux_io_enable)
  );
  ReadTableEntry ReadTable_0 ( // @[ReadMemoryController.scala 251:28]
    .clock(ReadTable_0_clock),
    .reset(ReadTable_0_reset),
    .io_NodeReq_ready(ReadTable_0_io_NodeReq_ready),
    .io_NodeReq_valid(ReadTable_0_io_NodeReq_valid),
    .io_NodeReq_bits_RouteID(ReadTable_0_io_NodeReq_bits_RouteID),
    .io_NodeReq_bits_address(ReadTable_0_io_NodeReq_bits_address),
    .io_NodeReq_bits_taskID(ReadTable_0_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(ReadTable_0_io_NodeReq_bits_Typ),
    .io_MemReq_ready(ReadTable_0_io_MemReq_ready),
    .io_MemReq_valid(ReadTable_0_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadTable_0_io_MemReq_bits_addr),
    .io_MemReq_bits_tag(ReadTable_0_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadTable_0_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadTable_0_io_MemReq_bits_iswrite),
    .io_MemResp_valid(ReadTable_0_io_MemResp_valid),
    .io_MemResp_data(ReadTable_0_io_MemResp_data),
    .io_output_ready(ReadTable_0_io_output_ready),
    .io_output_valid(ReadTable_0_io_output_valid),
    .io_output_bits_RouteID(ReadTable_0_io_output_bits_RouteID),
    .io_output_bits_data(ReadTable_0_io_output_bits_data),
    .io_free(ReadTable_0_io_free)
  );
  ReadTableEntry_1 ReadTable_1 ( // @[ReadMemoryController.scala 251:28]
    .clock(ReadTable_1_clock),
    .reset(ReadTable_1_reset),
    .io_NodeReq_ready(ReadTable_1_io_NodeReq_ready),
    .io_NodeReq_valid(ReadTable_1_io_NodeReq_valid),
    .io_NodeReq_bits_RouteID(ReadTable_1_io_NodeReq_bits_RouteID),
    .io_NodeReq_bits_address(ReadTable_1_io_NodeReq_bits_address),
    .io_NodeReq_bits_taskID(ReadTable_1_io_NodeReq_bits_taskID),
    .io_NodeReq_bits_Typ(ReadTable_1_io_NodeReq_bits_Typ),
    .io_MemReq_ready(ReadTable_1_io_MemReq_ready),
    .io_MemReq_valid(ReadTable_1_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadTable_1_io_MemReq_bits_addr),
    .io_MemReq_bits_tag(ReadTable_1_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadTable_1_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadTable_1_io_MemReq_bits_iswrite),
    .io_MemResp_valid(ReadTable_1_io_MemResp_valid),
    .io_MemResp_data(ReadTable_1_io_MemResp_data),
    .io_output_ready(ReadTable_1_io_output_ready),
    .io_output_valid(ReadTable_1_io_output_valid),
    .io_output_bits_RouteID(ReadTable_1_io_output_bits_RouteID),
    .io_output_bits_data(ReadTable_1_io_output_bits_data),
    .io_free(ReadTable_1_io_free)
  );
  assign io_ReadIn_0_ready = in_arb_io_in_0_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_1_ready = in_arb_io_in_1_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_2_ready = in_arb_io_in_2_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_3_ready = in_arb_io_in_3_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_4_ready = in_arb_io_in_4_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_5_ready = in_arb_io_in_5_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_6_ready = in_arb_io_in_6_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_7_ready = in_arb_io_in_7_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_8_ready = in_arb_io_in_8_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_9_ready = in_arb_io_in_9_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_10_ready = in_arb_io_in_10_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_11_ready = in_arb_io_in_11_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_12_ready = in_arb_io_in_12_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_13_ready = in_arb_io_in_13_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_14_ready = in_arb_io_in_14_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_15_ready = in_arb_io_in_15_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_16_ready = in_arb_io_in_16_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_17_ready = in_arb_io_in_17_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadIn_18_ready = in_arb_io_in_18_ready; // @[ReadMemoryController.scala 240:21]
  assign io_ReadOut_0_valid = out_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_0_data = out_demux_io_outputs_0_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_1_valid = out_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_1_data = out_demux_io_outputs_1_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_2_valid = out_demux_io_outputs_2_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_2_data = out_demux_io_outputs_2_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_3_valid = out_demux_io_outputs_3_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_3_data = out_demux_io_outputs_3_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_4_valid = out_demux_io_outputs_4_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_4_data = out_demux_io_outputs_4_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_5_valid = out_demux_io_outputs_5_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_5_data = out_demux_io_outputs_5_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_6_valid = out_demux_io_outputs_6_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_6_data = out_demux_io_outputs_6_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_7_valid = out_demux_io_outputs_7_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_7_data = out_demux_io_outputs_7_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_8_valid = out_demux_io_outputs_8_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_8_data = out_demux_io_outputs_8_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_9_valid = out_demux_io_outputs_9_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_9_data = out_demux_io_outputs_9_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_10_valid = out_demux_io_outputs_10_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_10_data = out_demux_io_outputs_10_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_11_valid = out_demux_io_outputs_11_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_11_data = out_demux_io_outputs_11_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_12_valid = out_demux_io_outputs_12_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_12_data = out_demux_io_outputs_12_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_13_valid = out_demux_io_outputs_13_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_13_data = out_demux_io_outputs_13_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_14_valid = out_demux_io_outputs_14_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_14_data = out_demux_io_outputs_14_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_15_valid = out_demux_io_outputs_15_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_15_data = out_demux_io_outputs_15_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_16_valid = out_demux_io_outputs_16_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_16_data = out_demux_io_outputs_16_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_17_valid = out_demux_io_outputs_17_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_17_data = out_demux_io_outputs_17_data; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_18_valid = out_demux_io_outputs_18_valid; // @[ReadMemoryController.scala 241:19]
  assign io_ReadOut_18_data = out_demux_io_outputs_18_data; // @[ReadMemoryController.scala 241:19]
  assign io_MemReq_valid = cachereq_arb_io_out_valid; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_addr = cachereq_arb_io_out_bits_addr; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_data = cachereq_arb_io_out_bits_data; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_mask = cachereq_arb_io_out_bits_mask; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_tag = cachereq_arb_io_out_bits_tag; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_taskID = cachereq_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 288:13]
  assign io_MemReq_bits_iswrite = cachereq_arb_io_out_bits_iswrite; // @[ReadMemoryController.scala 288:13]
  assign in_arb_clock = clock;
  assign in_arb_io_in_0_valid = io_ReadIn_0_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_0_bits_address = io_ReadIn_0_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_0_bits_taskID = io_ReadIn_0_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_1_valid = io_ReadIn_1_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_1_bits_address = io_ReadIn_1_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_1_bits_taskID = io_ReadIn_1_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_2_valid = io_ReadIn_2_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_2_bits_address = io_ReadIn_2_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_2_bits_taskID = io_ReadIn_2_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_3_valid = io_ReadIn_3_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_3_bits_address = io_ReadIn_3_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_3_bits_taskID = io_ReadIn_3_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_4_valid = io_ReadIn_4_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_4_bits_address = io_ReadIn_4_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_4_bits_taskID = io_ReadIn_4_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_5_valid = io_ReadIn_5_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_5_bits_address = io_ReadIn_5_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_5_bits_taskID = io_ReadIn_5_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_6_valid = io_ReadIn_6_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_6_bits_address = io_ReadIn_6_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_6_bits_taskID = io_ReadIn_6_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_7_valid = io_ReadIn_7_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_7_bits_address = io_ReadIn_7_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_7_bits_taskID = io_ReadIn_7_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_8_valid = io_ReadIn_8_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_8_bits_address = io_ReadIn_8_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_8_bits_taskID = io_ReadIn_8_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_9_valid = io_ReadIn_9_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_9_bits_address = io_ReadIn_9_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_9_bits_taskID = io_ReadIn_9_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_10_valid = io_ReadIn_10_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_10_bits_address = io_ReadIn_10_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_10_bits_taskID = io_ReadIn_10_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_11_valid = io_ReadIn_11_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_11_bits_address = io_ReadIn_11_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_11_bits_taskID = io_ReadIn_11_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_12_valid = io_ReadIn_12_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_12_bits_address = io_ReadIn_12_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_12_bits_taskID = io_ReadIn_12_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_13_valid = io_ReadIn_13_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_13_bits_address = io_ReadIn_13_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_13_bits_taskID = io_ReadIn_13_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_14_valid = io_ReadIn_14_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_14_bits_address = io_ReadIn_14_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_14_bits_taskID = io_ReadIn_14_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_15_valid = io_ReadIn_15_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_15_bits_address = io_ReadIn_15_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_15_bits_taskID = io_ReadIn_15_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_16_valid = io_ReadIn_16_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_16_bits_address = io_ReadIn_16_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_16_bits_taskID = io_ReadIn_16_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_17_valid = io_ReadIn_17_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_17_bits_address = io_ReadIn_17_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_17_bits_taskID = io_ReadIn_17_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_18_valid = io_ReadIn_18_valid; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_18_bits_address = io_ReadIn_18_bits_address; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_in_18_bits_taskID = io_ReadIn_18_bits_taskID; // @[ReadMemoryController.scala 240:21]
  assign in_arb_io_out_ready = alloc_arb_io_out_valid; // @[ReadMemoryController.scala 283:23]
  assign alloc_arb_io_in_0_valid = ReadTable_0_io_free; // @[ReadMemoryController.scala 254:30]
  assign alloc_arb_io_in_1_valid = ReadTable_1_io_free; // @[ReadMemoryController.scala 254:30]
  assign alloc_arb_io_out_ready = in_arb_io_out_valid; // @[ReadMemoryController.scala 284:26]
  assign cachereq_arb_io_in_0_valid = ReadTable_0_io_MemReq_valid; // @[ReadMemoryController.scala 260:33]
  assign cachereq_arb_io_in_0_bits_addr = ReadTable_0_io_MemReq_bits_addr; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_data = 32'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_mask = 4'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_tag = ReadTable_0_io_MemReq_bits_tag; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_taskID = ReadTable_0_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_0_bits_iswrite = ReadTable_0_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_valid = ReadTable_1_io_MemReq_valid; // @[ReadMemoryController.scala 260:33]
  assign cachereq_arb_io_in_1_bits_addr = ReadTable_1_io_MemReq_bits_addr; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_data = 32'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_mask = 4'h0; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_tag = ReadTable_1_io_MemReq_bits_tag; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_taskID = ReadTable_1_io_MemReq_bits_taskID; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_in_1_bits_iswrite = ReadTable_1_io_MemReq_bits_iswrite; // @[ReadMemoryController.scala 261:32]
  assign cachereq_arb_io_out_ready = io_MemReq_ready; // @[ReadMemoryController.scala 288:13]
  assign cacheresp_demux_io_en = io_MemResp_valid; // @[ReadMemoryController.scala 291:25]
  assign cacheresp_demux_io_input_data = io_MemResp_bits_data; // @[ReadMemoryController.scala 292:28]
  assign cacheresp_demux_io_input_tag = io_MemResp_bits_tag; // @[ReadMemoryController.scala 292:28]
  assign cacheresp_demux_io_sel = io_MemResp_bits_tag[0]; // @[ReadMemoryController.scala 293:26]
  assign out_arb_clock = clock;
  assign out_arb_io_in_0_valid = ReadTable_0_io_output_valid; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_0_bits_RouteID = ReadTable_0_io_output_bits_RouteID; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_0_bits_data = ReadTable_0_io_output_bits_data; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_1_valid = ReadTable_1_io_output_valid; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_1_bits_RouteID = ReadTable_1_io_output_bits_RouteID; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_in_1_bits_data = ReadTable_1_io_output_bits_data; // @[ReadMemoryController.scala 268:22]
  assign out_arb_io_out_ready = 1'h1; // @[ReadMemoryController.scala 296:24]
  assign out_demux_clock = clock;
  assign out_demux_reset = reset;
  assign out_demux_io_input_RouteID = out_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 298:22]
  assign out_demux_io_input_data = out_arb_io_out_bits_data; // @[ReadMemoryController.scala 298:22]
  assign out_demux_io_enable = out_arb_io_out_ready & out_arb_io_out_valid; // @[ReadMemoryController.scala 297:23]
  assign ReadTable_0_clock = clock;
  assign ReadTable_0_reset = reset;
  assign ReadTable_0_io_NodeReq_valid = alloc_arb_io_in_0_ready & alloc_arb_io_in_0_valid; // @[ReadMemoryController.scala 256:33]
  assign ReadTable_0_io_NodeReq_bits_RouteID = in_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_0_io_MemReq_ready = cachereq_arb_io_in_0_ready; // @[ReadMemoryController.scala 262:32]
  assign ReadTable_0_io_MemResp_valid = cacheresp_demux_io_outputs_0_valid; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_0_io_MemResp_data = cacheresp_demux_io_outputs_0_data; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_0_io_output_ready = out_arb_io_in_0_ready; // @[ReadMemoryController.scala 268:22]
  assign ReadTable_1_clock = clock;
  assign ReadTable_1_reset = reset;
  assign ReadTable_1_io_NodeReq_valid = alloc_arb_io_in_1_ready & alloc_arb_io_in_1_valid; // @[ReadMemoryController.scala 256:33]
  assign ReadTable_1_io_NodeReq_bits_RouteID = in_arb_io_out_bits_RouteID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_NodeReq_bits_address = in_arb_io_out_bits_address; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_NodeReq_bits_taskID = in_arb_io_out_bits_taskID; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_NodeReq_bits_Typ = in_arb_io_out_bits_Typ; // @[ReadMemoryController.scala 257:32]
  assign ReadTable_1_io_MemReq_ready = cachereq_arb_io_in_1_ready; // @[ReadMemoryController.scala 262:32]
  assign ReadTable_1_io_MemResp_valid = cacheresp_demux_io_outputs_1_valid; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_1_io_MemResp_data = cacheresp_demux_io_outputs_1_data; // @[ReadMemoryController.scala 265:27]
  assign ReadTable_1_io_output_ready = out_arb_io_in_1_ready; // @[ReadMemoryController.scala 268:22]
endmodule
module RRArbiter_2(
  input         clock,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [31:0] io_in_0_bits_data,
  input  [3:0]  io_in_0_bits_mask,
  input  [7:0]  io_in_0_bits_tag,
  input  [4:0]  io_in_0_bits_taskID,
  input         io_in_0_bits_iswrite,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [31:0] io_in_1_bits_data,
  input  [3:0]  io_in_1_bits_mask,
  input  [7:0]  io_in_1_bits_tag,
  input  [4:0]  io_in_1_bits_taskID,
  input         io_in_1_bits_iswrite,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [31:0] io_out_bits_data,
  output [3:0]  io_out_bits_mask,
  output [7:0]  io_out_bits_tag,
  output [4:0]  io_out_bits_taskID,
  output        io_out_bits_iswrite,
  output        io_chosen
);
  wire  _T; // @[Decoupled.scala 40:37]
  reg  _T_1; // @[Reg.scala 15:16]
  reg [31:0] _RAND_0;
  wire  _T_3; // @[Arbiter.scala 67:57]
  wire  _T_5; // @[Arbiter.scala 68:83]
  wire  _T_7; // @[Arbiter.scala 31:68]
  wire  _T_9; // @[Arbiter.scala 31:78]
  wire  _T_10; // @[Arbiter.scala 31:78]
  wire  _T_14; // @[Arbiter.scala 72:50]
  wire  _GEN_19; // @[Arbiter.scala 77:27]
  assign _T = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = 1'h1 > _T_1; // @[Arbiter.scala 67:57]
  assign _T_5 = io_in_1_valid & _T_3; // @[Arbiter.scala 68:83]
  assign _T_7 = _T_5 | io_in_0_valid; // @[Arbiter.scala 31:68]
  assign _T_9 = _T_5 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_10 = _T_7 == 1'h0; // @[Arbiter.scala 31:78]
  assign _T_14 = _T_3 | _T_10; // @[Arbiter.scala 72:50]
  assign _GEN_19 = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 77:27]
  assign io_in_0_ready = _T_9 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_in_1_ready = _T_14 & io_out_ready; // @[Arbiter.scala 60:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15]
  assign io_out_bits_data = io_chosen ? io_in_1_bits_data : io_in_0_bits_data; // @[Arbiter.scala 42:15]
  assign io_out_bits_mask = io_chosen ? io_in_1_bits_mask : io_in_0_bits_mask; // @[Arbiter.scala 42:15]
  assign io_out_bits_tag = io_chosen ? io_in_1_bits_tag : io_in_0_bits_tag; // @[Arbiter.scala 42:15]
  assign io_out_bits_taskID = io_chosen ? io_in_1_bits_taskID : io_in_0_bits_taskID; // @[Arbiter.scala 42:15]
  assign io_out_bits_iswrite = io_chosen ? io_in_1_bits_iswrite : io_in_0_bits_iswrite; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_5 | _GEN_19; // @[Arbiter.scala 40:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (_T) begin
      _T_1 <= io_chosen;
    end
  end
endmodule
module ReadWriteArbiter(
  input         clock,
  output        io_ReadMemReq_ready,
  input         io_ReadMemReq_valid,
  input  [31:0] io_ReadMemReq_bits_addr,
  input  [31:0] io_ReadMemReq_bits_data,
  input  [3:0]  io_ReadMemReq_bits_mask,
  input  [7:0]  io_ReadMemReq_bits_tag,
  input  [4:0]  io_ReadMemReq_bits_taskID,
  input         io_ReadMemReq_bits_iswrite,
  output        io_WriteMemReq_ready,
  input         io_WriteMemReq_valid,
  input  [31:0] io_WriteMemReq_bits_addr,
  input  [31:0] io_WriteMemReq_bits_data,
  input  [3:0]  io_WriteMemReq_bits_mask,
  input  [7:0]  io_WriteMemReq_bits_tag,
  input  [4:0]  io_WriteMemReq_bits_taskID,
  input         io_WriteMemReq_bits_iswrite,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemResp_bits_iswrite,
  output        io_ReadMemResp_valid,
  output [31:0] io_ReadMemResp_bits_data,
  output [7:0]  io_ReadMemResp_bits_tag,
  output        io_WriteMemResp_valid,
  output [31:0] io_WriteMemResp_bits_data,
  output [7:0]  io_WriteMemResp_bits_tag,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite
);
  wire  cachereq_arb_clock; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_0_ready; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_0_valid; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_0_bits_addr; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_0_bits_data; // @[ReadWriteArbiter.scala 48:31]
  wire [3:0] cachereq_arb_io_in_0_bits_mask; // @[ReadWriteArbiter.scala 48:31]
  wire [7:0] cachereq_arb_io_in_0_bits_tag; // @[ReadWriteArbiter.scala 48:31]
  wire [4:0] cachereq_arb_io_in_0_bits_taskID; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_0_bits_iswrite; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_1_ready; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_1_valid; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_1_bits_addr; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_in_1_bits_data; // @[ReadWriteArbiter.scala 48:31]
  wire [3:0] cachereq_arb_io_in_1_bits_mask; // @[ReadWriteArbiter.scala 48:31]
  wire [7:0] cachereq_arb_io_in_1_bits_tag; // @[ReadWriteArbiter.scala 48:31]
  wire [4:0] cachereq_arb_io_in_1_bits_taskID; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_in_1_bits_iswrite; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_out_ready; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_out_valid; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_out_bits_addr; // @[ReadWriteArbiter.scala 48:31]
  wire [31:0] cachereq_arb_io_out_bits_data; // @[ReadWriteArbiter.scala 48:31]
  wire [3:0] cachereq_arb_io_out_bits_mask; // @[ReadWriteArbiter.scala 48:31]
  wire [7:0] cachereq_arb_io_out_bits_tag; // @[ReadWriteArbiter.scala 48:31]
  wire [4:0] cachereq_arb_io_out_bits_taskID; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_out_bits_iswrite; // @[ReadWriteArbiter.scala 48:31]
  wire  cachereq_arb_io_chosen; // @[ReadWriteArbiter.scala 48:31]
  wire  cacheresp_demux_io_en; // @[ReadWriteArbiter.scala 50:31]
  wire [31:0] cacheresp_demux_io_input_data; // @[ReadWriteArbiter.scala 50:31]
  wire [7:0] cacheresp_demux_io_input_tag; // @[ReadWriteArbiter.scala 50:31]
  wire  cacheresp_demux_io_sel; // @[ReadWriteArbiter.scala 50:31]
  wire  cacheresp_demux_io_outputs_0_valid; // @[ReadWriteArbiter.scala 50:31]
  wire [31:0] cacheresp_demux_io_outputs_0_data; // @[ReadWriteArbiter.scala 50:31]
  wire [7:0] cacheresp_demux_io_outputs_0_tag; // @[ReadWriteArbiter.scala 50:31]
  wire  cacheresp_demux_io_outputs_1_valid; // @[ReadWriteArbiter.scala 50:31]
  wire [31:0] cacheresp_demux_io_outputs_1_data; // @[ReadWriteArbiter.scala 50:31]
  wire [7:0] cacheresp_demux_io_outputs_1_tag; // @[ReadWriteArbiter.scala 50:31]
  RRArbiter_2 cachereq_arb ( // @[ReadWriteArbiter.scala 48:31]
    .clock(cachereq_arb_clock),
    .io_in_0_ready(cachereq_arb_io_in_0_ready),
    .io_in_0_valid(cachereq_arb_io_in_0_valid),
    .io_in_0_bits_addr(cachereq_arb_io_in_0_bits_addr),
    .io_in_0_bits_data(cachereq_arb_io_in_0_bits_data),
    .io_in_0_bits_mask(cachereq_arb_io_in_0_bits_mask),
    .io_in_0_bits_tag(cachereq_arb_io_in_0_bits_tag),
    .io_in_0_bits_taskID(cachereq_arb_io_in_0_bits_taskID),
    .io_in_0_bits_iswrite(cachereq_arb_io_in_0_bits_iswrite),
    .io_in_1_ready(cachereq_arb_io_in_1_ready),
    .io_in_1_valid(cachereq_arb_io_in_1_valid),
    .io_in_1_bits_addr(cachereq_arb_io_in_1_bits_addr),
    .io_in_1_bits_data(cachereq_arb_io_in_1_bits_data),
    .io_in_1_bits_mask(cachereq_arb_io_in_1_bits_mask),
    .io_in_1_bits_tag(cachereq_arb_io_in_1_bits_tag),
    .io_in_1_bits_taskID(cachereq_arb_io_in_1_bits_taskID),
    .io_in_1_bits_iswrite(cachereq_arb_io_in_1_bits_iswrite),
    .io_out_ready(cachereq_arb_io_out_ready),
    .io_out_valid(cachereq_arb_io_out_valid),
    .io_out_bits_addr(cachereq_arb_io_out_bits_addr),
    .io_out_bits_data(cachereq_arb_io_out_bits_data),
    .io_out_bits_mask(cachereq_arb_io_out_bits_mask),
    .io_out_bits_tag(cachereq_arb_io_out_bits_tag),
    .io_out_bits_taskID(cachereq_arb_io_out_bits_taskID),
    .io_out_bits_iswrite(cachereq_arb_io_out_bits_iswrite),
    .io_chosen(cachereq_arb_io_chosen)
  );
  Demux cacheresp_demux ( // @[ReadWriteArbiter.scala 50:31]
    .io_en(cacheresp_demux_io_en),
    .io_input_data(cacheresp_demux_io_input_data),
    .io_input_tag(cacheresp_demux_io_input_tag),
    .io_sel(cacheresp_demux_io_sel),
    .io_outputs_0_valid(cacheresp_demux_io_outputs_0_valid),
    .io_outputs_0_data(cacheresp_demux_io_outputs_0_data),
    .io_outputs_0_tag(cacheresp_demux_io_outputs_0_tag),
    .io_outputs_1_valid(cacheresp_demux_io_outputs_1_valid),
    .io_outputs_1_data(cacheresp_demux_io_outputs_1_data),
    .io_outputs_1_tag(cacheresp_demux_io_outputs_1_tag)
  );
  assign io_ReadMemReq_ready = cachereq_arb_io_in_0_ready; // @[ReadWriteArbiter.scala 57:29]
  assign io_WriteMemReq_ready = cachereq_arb_io_in_1_ready; // @[ReadWriteArbiter.scala 58:29]
  assign io_ReadMemResp_valid = cacheresp_demux_io_outputs_0_valid; // @[ReadWriteArbiter.scala 69:24]
  assign io_ReadMemResp_bits_data = cacheresp_demux_io_outputs_0_data; // @[ReadWriteArbiter.scala 68:23]
  assign io_ReadMemResp_bits_tag = cacheresp_demux_io_outputs_0_tag; // @[ReadWriteArbiter.scala 68:23]
  assign io_WriteMemResp_valid = cacheresp_demux_io_outputs_1_valid; // @[ReadWriteArbiter.scala 71:25]
  assign io_WriteMemResp_bits_data = cacheresp_demux_io_outputs_1_data; // @[ReadWriteArbiter.scala 70:24]
  assign io_WriteMemResp_bits_tag = cacheresp_demux_io_outputs_1_tag; // @[ReadWriteArbiter.scala 70:24]
  assign io_MemReq_valid = cachereq_arb_io_out_valid; // @[ReadWriteArbiter.scala 62:19]
  assign io_MemReq_bits_addr = cachereq_arb_io_out_bits_addr; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_data = cachereq_arb_io_out_bits_data; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_mask = cachereq_arb_io_out_bits_mask; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_tag = cachereq_arb_io_out_bits_tag; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_taskID = cachereq_arb_io_out_bits_taskID; // @[ReadWriteArbiter.scala 61:18]
  assign io_MemReq_bits_iswrite = cachereq_arb_io_out_bits_iswrite; // @[ReadWriteArbiter.scala 61:18]
  assign cachereq_arb_clock = clock;
  assign cachereq_arb_io_in_0_valid = io_ReadMemReq_valid; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_addr = io_ReadMemReq_bits_addr; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_data = io_ReadMemReq_bits_data; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_mask = io_ReadMemReq_bits_mask; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_tag = io_ReadMemReq_bits_tag; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_taskID = io_ReadMemReq_bits_taskID; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_0_bits_iswrite = io_ReadMemReq_bits_iswrite; // @[ReadWriteArbiter.scala 57:29]
  assign cachereq_arb_io_in_1_valid = io_WriteMemReq_valid; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_addr = io_WriteMemReq_bits_addr; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_data = io_WriteMemReq_bits_data; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_mask = io_WriteMemReq_bits_mask; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_tag = io_WriteMemReq_bits_tag; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_taskID = io_WriteMemReq_bits_taskID; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_in_1_bits_iswrite = io_WriteMemReq_bits_iswrite; // @[ReadWriteArbiter.scala 58:29]
  assign cachereq_arb_io_out_ready = io_MemReq_ready; // @[ReadWriteArbiter.scala 60:29]
  assign cacheresp_demux_io_en = io_MemResp_valid; // @[ReadWriteArbiter.scala 76:25]
  assign cacheresp_demux_io_input_data = io_MemResp_bits_data; // @[ReadWriteArbiter.scala 77:28]
  assign cacheresp_demux_io_input_tag = io_MemResp_bits_tag; // @[ReadWriteArbiter.scala 77:28]
  assign cacheresp_demux_io_sel = io_MemResp_bits_iswrite; // @[ReadWriteArbiter.scala 80:26]
endmodule
module UnifiedController(
  input         clock,
  input         reset,
  output        io_WriteIn_0_ready,
  input         io_WriteIn_0_valid,
  input  [21:0] io_WriteIn_0_bits_address,
  input  [31:0] io_WriteIn_0_bits_data,
  input  [4:0]  io_WriteIn_0_bits_taskID,
  output        io_WriteIn_1_ready,
  input         io_WriteIn_1_valid,
  input  [21:0] io_WriteIn_1_bits_address,
  input  [31:0] io_WriteIn_1_bits_data,
  input  [4:0]  io_WriteIn_1_bits_taskID,
  output        io_WriteIn_2_ready,
  input         io_WriteIn_2_valid,
  input  [21:0] io_WriteIn_2_bits_address,
  input  [31:0] io_WriteIn_2_bits_data,
  input  [4:0]  io_WriteIn_2_bits_taskID,
  output        io_WriteIn_3_ready,
  input         io_WriteIn_3_valid,
  input  [21:0] io_WriteIn_3_bits_address,
  input  [31:0] io_WriteIn_3_bits_data,
  input  [4:0]  io_WriteIn_3_bits_taskID,
  output        io_WriteIn_4_ready,
  input         io_WriteIn_4_valid,
  input  [21:0] io_WriteIn_4_bits_address,
  input  [31:0] io_WriteIn_4_bits_data,
  input  [4:0]  io_WriteIn_4_bits_taskID,
  output        io_WriteIn_5_ready,
  input         io_WriteIn_5_valid,
  input  [21:0] io_WriteIn_5_bits_address,
  input  [31:0] io_WriteIn_5_bits_data,
  input  [4:0]  io_WriteIn_5_bits_taskID,
  output        io_WriteIn_6_ready,
  input         io_WriteIn_6_valid,
  input  [21:0] io_WriteIn_6_bits_address,
  input  [31:0] io_WriteIn_6_bits_data,
  input  [4:0]  io_WriteIn_6_bits_taskID,
  output        io_WriteIn_7_ready,
  input         io_WriteIn_7_valid,
  input  [21:0] io_WriteIn_7_bits_address,
  input  [31:0] io_WriteIn_7_bits_data,
  input  [4:0]  io_WriteIn_7_bits_taskID,
  output        io_WriteIn_8_ready,
  input         io_WriteIn_8_valid,
  input  [21:0] io_WriteIn_8_bits_address,
  input  [31:0] io_WriteIn_8_bits_data,
  input  [4:0]  io_WriteIn_8_bits_taskID,
  output        io_WriteOut_0_valid,
  output        io_WriteOut_1_valid,
  output        io_WriteOut_2_valid,
  output        io_WriteOut_3_valid,
  output        io_WriteOut_4_valid,
  output        io_WriteOut_5_valid,
  output        io_WriteOut_6_valid,
  output        io_WriteOut_7_valid,
  output        io_WriteOut_8_valid,
  output        io_ReadIn_0_ready,
  input         io_ReadIn_0_valid,
  input  [31:0] io_ReadIn_0_bits_address,
  input  [4:0]  io_ReadIn_0_bits_taskID,
  output        io_ReadIn_1_ready,
  input         io_ReadIn_1_valid,
  input  [31:0] io_ReadIn_1_bits_address,
  input  [4:0]  io_ReadIn_1_bits_taskID,
  output        io_ReadIn_2_ready,
  input         io_ReadIn_2_valid,
  input  [31:0] io_ReadIn_2_bits_address,
  input  [4:0]  io_ReadIn_2_bits_taskID,
  output        io_ReadIn_3_ready,
  input         io_ReadIn_3_valid,
  input  [31:0] io_ReadIn_3_bits_address,
  input  [4:0]  io_ReadIn_3_bits_taskID,
  output        io_ReadIn_4_ready,
  input         io_ReadIn_4_valid,
  input  [31:0] io_ReadIn_4_bits_address,
  input  [4:0]  io_ReadIn_4_bits_taskID,
  output        io_ReadIn_5_ready,
  input         io_ReadIn_5_valid,
  input  [31:0] io_ReadIn_5_bits_address,
  input  [4:0]  io_ReadIn_5_bits_taskID,
  output        io_ReadIn_6_ready,
  input         io_ReadIn_6_valid,
  input  [31:0] io_ReadIn_6_bits_address,
  input  [4:0]  io_ReadIn_6_bits_taskID,
  output        io_ReadIn_7_ready,
  input         io_ReadIn_7_valid,
  input  [31:0] io_ReadIn_7_bits_address,
  input  [4:0]  io_ReadIn_7_bits_taskID,
  output        io_ReadIn_8_ready,
  input         io_ReadIn_8_valid,
  input  [31:0] io_ReadIn_8_bits_address,
  input  [4:0]  io_ReadIn_8_bits_taskID,
  output        io_ReadIn_9_ready,
  input         io_ReadIn_9_valid,
  input  [31:0] io_ReadIn_9_bits_address,
  input  [4:0]  io_ReadIn_9_bits_taskID,
  output        io_ReadIn_10_ready,
  input         io_ReadIn_10_valid,
  input  [31:0] io_ReadIn_10_bits_address,
  input  [4:0]  io_ReadIn_10_bits_taskID,
  output        io_ReadIn_11_ready,
  input         io_ReadIn_11_valid,
  input  [31:0] io_ReadIn_11_bits_address,
  input  [4:0]  io_ReadIn_11_bits_taskID,
  output        io_ReadIn_12_ready,
  input         io_ReadIn_12_valid,
  input  [31:0] io_ReadIn_12_bits_address,
  input  [4:0]  io_ReadIn_12_bits_taskID,
  output        io_ReadIn_13_ready,
  input         io_ReadIn_13_valid,
  input  [31:0] io_ReadIn_13_bits_address,
  input  [4:0]  io_ReadIn_13_bits_taskID,
  output        io_ReadIn_14_ready,
  input         io_ReadIn_14_valid,
  input  [31:0] io_ReadIn_14_bits_address,
  input  [4:0]  io_ReadIn_14_bits_taskID,
  output        io_ReadIn_15_ready,
  input         io_ReadIn_15_valid,
  input  [31:0] io_ReadIn_15_bits_address,
  input  [4:0]  io_ReadIn_15_bits_taskID,
  output        io_ReadIn_16_ready,
  input         io_ReadIn_16_valid,
  input  [31:0] io_ReadIn_16_bits_address,
  input  [4:0]  io_ReadIn_16_bits_taskID,
  output        io_ReadIn_17_ready,
  input         io_ReadIn_17_valid,
  input  [31:0] io_ReadIn_17_bits_address,
  input  [4:0]  io_ReadIn_17_bits_taskID,
  output        io_ReadIn_18_ready,
  input         io_ReadIn_18_valid,
  input  [31:0] io_ReadIn_18_bits_address,
  input  [4:0]  io_ReadIn_18_bits_taskID,
  output        io_ReadOut_0_valid,
  output [31:0] io_ReadOut_0_data,
  output        io_ReadOut_1_valid,
  output [31:0] io_ReadOut_1_data,
  output        io_ReadOut_2_valid,
  output [31:0] io_ReadOut_2_data,
  output        io_ReadOut_3_valid,
  output [31:0] io_ReadOut_3_data,
  output        io_ReadOut_4_valid,
  output [31:0] io_ReadOut_4_data,
  output        io_ReadOut_5_valid,
  output [31:0] io_ReadOut_5_data,
  output        io_ReadOut_6_valid,
  output [31:0] io_ReadOut_6_data,
  output        io_ReadOut_7_valid,
  output [31:0] io_ReadOut_7_data,
  output        io_ReadOut_8_valid,
  output [31:0] io_ReadOut_8_data,
  output        io_ReadOut_9_valid,
  output [31:0] io_ReadOut_9_data,
  output        io_ReadOut_10_valid,
  output [31:0] io_ReadOut_10_data,
  output        io_ReadOut_11_valid,
  output [31:0] io_ReadOut_11_data,
  output        io_ReadOut_12_valid,
  output [31:0] io_ReadOut_12_data,
  output        io_ReadOut_13_valid,
  output [31:0] io_ReadOut_13_data,
  output        io_ReadOut_14_valid,
  output [31:0] io_ReadOut_14_data,
  output        io_ReadOut_15_valid,
  output [31:0] io_ReadOut_15_data,
  output        io_ReadOut_16_valid,
  output [31:0] io_ReadOut_16_data,
  output        io_ReadOut_17_valid,
  output [31:0] io_ReadOut_17_data,
  output        io_ReadOut_18_valid,
  output [31:0] io_ReadOut_18_data,
  input         io_MemResp_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemResp_bits_iswrite,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite
);
  wire  WriteController_clock; // @[UnifiedController.scala 53:32]
  wire  WriteController_reset; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_0_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_0_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_0_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_0_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_0_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_1_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_1_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_1_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_1_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_1_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_2_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_2_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_2_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_2_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_2_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_3_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_3_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_3_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_3_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_3_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_4_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_4_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_4_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_4_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_4_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_5_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_5_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_5_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_5_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_5_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_6_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_6_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_6_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_6_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_6_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_7_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_7_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_7_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_7_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_7_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_8_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteIn_8_valid; // @[UnifiedController.scala 53:32]
  wire [21:0] WriteController_io_WriteIn_8_bits_address; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_WriteIn_8_bits_data; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_WriteIn_8_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_0_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_1_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_2_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_3_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_4_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_5_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_6_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_7_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_WriteOut_8_valid; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_MemReq_ready; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_MemReq_valid; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_MemReq_bits_addr; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_MemReq_bits_data; // @[UnifiedController.scala 53:32]
  wire [3:0] WriteController_io_MemReq_bits_mask; // @[UnifiedController.scala 53:32]
  wire [7:0] WriteController_io_MemReq_bits_tag; // @[UnifiedController.scala 53:32]
  wire [4:0] WriteController_io_MemReq_bits_taskID; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 53:32]
  wire  WriteController_io_MemResp_valid; // @[UnifiedController.scala 53:32]
  wire [31:0] WriteController_io_MemResp_bits_data; // @[UnifiedController.scala 53:32]
  wire [7:0] WriteController_io_MemResp_bits_tag; // @[UnifiedController.scala 53:32]
  wire  ReadController_clock; // @[UnifiedController.scala 54:32]
  wire  ReadController_reset; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_0_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_0_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_0_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_0_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_1_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_1_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_1_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_1_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_2_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_2_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_2_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_2_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_3_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_3_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_3_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_3_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_4_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_4_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_4_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_4_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_5_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_5_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_5_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_5_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_6_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_6_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_6_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_6_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_7_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_7_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_7_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_7_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_8_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_8_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_8_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_8_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_9_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_9_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_9_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_9_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_10_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_10_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_10_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_10_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_11_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_11_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_11_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_11_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_12_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_12_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_12_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_12_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_13_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_13_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_13_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_13_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_14_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_14_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_14_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_14_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_15_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_15_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_15_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_15_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_16_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_16_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_16_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_16_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_17_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_17_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_17_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_17_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_18_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadIn_18_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadIn_18_bits_address; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_ReadIn_18_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_0_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_0_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_1_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_1_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_2_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_2_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_3_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_3_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_4_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_4_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_5_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_5_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_6_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_6_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_7_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_7_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_8_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_8_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_9_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_9_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_10_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_10_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_11_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_11_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_12_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_12_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_13_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_13_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_14_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_14_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_15_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_15_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_16_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_16_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_17_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_17_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_ReadOut_18_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_ReadOut_18_data; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_MemReq_ready; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_MemReq_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_MemReq_bits_addr; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_MemReq_bits_data; // @[UnifiedController.scala 54:32]
  wire [3:0] ReadController_io_MemReq_bits_mask; // @[UnifiedController.scala 54:32]
  wire [7:0] ReadController_io_MemReq_bits_tag; // @[UnifiedController.scala 54:32]
  wire [4:0] ReadController_io_MemReq_bits_taskID; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 54:32]
  wire  ReadController_io_MemResp_valid; // @[UnifiedController.scala 54:32]
  wire [31:0] ReadController_io_MemResp_bits_data; // @[UnifiedController.scala 54:32]
  wire [7:0] ReadController_io_MemResp_bits_tag; // @[UnifiedController.scala 54:32]
  wire  ReadWriteArbiter_clock; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_ReadMemReq_ready; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_ReadMemReq_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_ReadMemReq_bits_addr; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_ReadMemReq_bits_data; // @[UnifiedController.scala 55:32]
  wire [3:0] ReadWriteArbiter_io_ReadMemReq_bits_mask; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_ReadMemReq_bits_tag; // @[UnifiedController.scala 55:32]
  wire [4:0] ReadWriteArbiter_io_ReadMemReq_bits_taskID; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_ReadMemReq_bits_iswrite; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_WriteMemReq_ready; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_WriteMemReq_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_WriteMemReq_bits_addr; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_WriteMemReq_bits_data; // @[UnifiedController.scala 55:32]
  wire [3:0] ReadWriteArbiter_io_WriteMemReq_bits_mask; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_WriteMemReq_bits_tag; // @[UnifiedController.scala 55:32]
  wire [4:0] ReadWriteArbiter_io_WriteMemReq_bits_taskID; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_WriteMemReq_bits_iswrite; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemResp_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_MemResp_bits_data; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_MemResp_bits_tag; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemResp_bits_iswrite; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_ReadMemResp_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_ReadMemResp_bits_data; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_ReadMemResp_bits_tag; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_WriteMemResp_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_WriteMemResp_bits_data; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_WriteMemResp_bits_tag; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemReq_ready; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemReq_valid; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_MemReq_bits_addr; // @[UnifiedController.scala 55:32]
  wire [31:0] ReadWriteArbiter_io_MemReq_bits_data; // @[UnifiedController.scala 55:32]
  wire [3:0] ReadWriteArbiter_io_MemReq_bits_mask; // @[UnifiedController.scala 55:32]
  wire [7:0] ReadWriteArbiter_io_MemReq_bits_tag; // @[UnifiedController.scala 55:32]
  wire [4:0] ReadWriteArbiter_io_MemReq_bits_taskID; // @[UnifiedController.scala 55:32]
  wire  ReadWriteArbiter_io_MemReq_bits_iswrite; // @[UnifiedController.scala 55:32]
  wire  _T; // @[Decoupled.scala 40:37]
  wire  _T_1; // @[UnifiedController.scala 92:15]
  wire  _T_2; // @[UnifiedController.scala 92:15]
  wire  _GEN_0; // @[UnifiedController.scala 92:15]
  wire  _GEN_1; // @[UnifiedController.scala 94:15]
  wire  _GEN_2; // @[UnifiedController.scala 94:15]
  wire  _GEN_3; // @[UnifiedController.scala 100:15]
  wire  _GEN_4; // @[UnifiedController.scala 102:15]
  wire  _GEN_5; // @[UnifiedController.scala 102:15]
  WriteMemoryController WriteController ( // @[UnifiedController.scala 53:32]
    .clock(WriteController_clock),
    .reset(WriteController_reset),
    .io_WriteIn_0_ready(WriteController_io_WriteIn_0_ready),
    .io_WriteIn_0_valid(WriteController_io_WriteIn_0_valid),
    .io_WriteIn_0_bits_address(WriteController_io_WriteIn_0_bits_address),
    .io_WriteIn_0_bits_data(WriteController_io_WriteIn_0_bits_data),
    .io_WriteIn_0_bits_taskID(WriteController_io_WriteIn_0_bits_taskID),
    .io_WriteIn_1_ready(WriteController_io_WriteIn_1_ready),
    .io_WriteIn_1_valid(WriteController_io_WriteIn_1_valid),
    .io_WriteIn_1_bits_address(WriteController_io_WriteIn_1_bits_address),
    .io_WriteIn_1_bits_data(WriteController_io_WriteIn_1_bits_data),
    .io_WriteIn_1_bits_taskID(WriteController_io_WriteIn_1_bits_taskID),
    .io_WriteIn_2_ready(WriteController_io_WriteIn_2_ready),
    .io_WriteIn_2_valid(WriteController_io_WriteIn_2_valid),
    .io_WriteIn_2_bits_address(WriteController_io_WriteIn_2_bits_address),
    .io_WriteIn_2_bits_data(WriteController_io_WriteIn_2_bits_data),
    .io_WriteIn_2_bits_taskID(WriteController_io_WriteIn_2_bits_taskID),
    .io_WriteIn_3_ready(WriteController_io_WriteIn_3_ready),
    .io_WriteIn_3_valid(WriteController_io_WriteIn_3_valid),
    .io_WriteIn_3_bits_address(WriteController_io_WriteIn_3_bits_address),
    .io_WriteIn_3_bits_data(WriteController_io_WriteIn_3_bits_data),
    .io_WriteIn_3_bits_taskID(WriteController_io_WriteIn_3_bits_taskID),
    .io_WriteIn_4_ready(WriteController_io_WriteIn_4_ready),
    .io_WriteIn_4_valid(WriteController_io_WriteIn_4_valid),
    .io_WriteIn_4_bits_address(WriteController_io_WriteIn_4_bits_address),
    .io_WriteIn_4_bits_data(WriteController_io_WriteIn_4_bits_data),
    .io_WriteIn_4_bits_taskID(WriteController_io_WriteIn_4_bits_taskID),
    .io_WriteIn_5_ready(WriteController_io_WriteIn_5_ready),
    .io_WriteIn_5_valid(WriteController_io_WriteIn_5_valid),
    .io_WriteIn_5_bits_address(WriteController_io_WriteIn_5_bits_address),
    .io_WriteIn_5_bits_data(WriteController_io_WriteIn_5_bits_data),
    .io_WriteIn_5_bits_taskID(WriteController_io_WriteIn_5_bits_taskID),
    .io_WriteIn_6_ready(WriteController_io_WriteIn_6_ready),
    .io_WriteIn_6_valid(WriteController_io_WriteIn_6_valid),
    .io_WriteIn_6_bits_address(WriteController_io_WriteIn_6_bits_address),
    .io_WriteIn_6_bits_data(WriteController_io_WriteIn_6_bits_data),
    .io_WriteIn_6_bits_taskID(WriteController_io_WriteIn_6_bits_taskID),
    .io_WriteIn_7_ready(WriteController_io_WriteIn_7_ready),
    .io_WriteIn_7_valid(WriteController_io_WriteIn_7_valid),
    .io_WriteIn_7_bits_address(WriteController_io_WriteIn_7_bits_address),
    .io_WriteIn_7_bits_data(WriteController_io_WriteIn_7_bits_data),
    .io_WriteIn_7_bits_taskID(WriteController_io_WriteIn_7_bits_taskID),
    .io_WriteIn_8_ready(WriteController_io_WriteIn_8_ready),
    .io_WriteIn_8_valid(WriteController_io_WriteIn_8_valid),
    .io_WriteIn_8_bits_address(WriteController_io_WriteIn_8_bits_address),
    .io_WriteIn_8_bits_data(WriteController_io_WriteIn_8_bits_data),
    .io_WriteIn_8_bits_taskID(WriteController_io_WriteIn_8_bits_taskID),
    .io_WriteOut_0_valid(WriteController_io_WriteOut_0_valid),
    .io_WriteOut_1_valid(WriteController_io_WriteOut_1_valid),
    .io_WriteOut_2_valid(WriteController_io_WriteOut_2_valid),
    .io_WriteOut_3_valid(WriteController_io_WriteOut_3_valid),
    .io_WriteOut_4_valid(WriteController_io_WriteOut_4_valid),
    .io_WriteOut_5_valid(WriteController_io_WriteOut_5_valid),
    .io_WriteOut_6_valid(WriteController_io_WriteOut_6_valid),
    .io_WriteOut_7_valid(WriteController_io_WriteOut_7_valid),
    .io_WriteOut_8_valid(WriteController_io_WriteOut_8_valid),
    .io_MemReq_ready(WriteController_io_MemReq_ready),
    .io_MemReq_valid(WriteController_io_MemReq_valid),
    .io_MemReq_bits_addr(WriteController_io_MemReq_bits_addr),
    .io_MemReq_bits_data(WriteController_io_MemReq_bits_data),
    .io_MemReq_bits_mask(WriteController_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(WriteController_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(WriteController_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(WriteController_io_MemReq_bits_iswrite),
    .io_MemResp_valid(WriteController_io_MemResp_valid),
    .io_MemResp_bits_data(WriteController_io_MemResp_bits_data),
    .io_MemResp_bits_tag(WriteController_io_MemResp_bits_tag)
  );
  ReadMemoryController ReadController ( // @[UnifiedController.scala 54:32]
    .clock(ReadController_clock),
    .reset(ReadController_reset),
    .io_ReadIn_0_ready(ReadController_io_ReadIn_0_ready),
    .io_ReadIn_0_valid(ReadController_io_ReadIn_0_valid),
    .io_ReadIn_0_bits_address(ReadController_io_ReadIn_0_bits_address),
    .io_ReadIn_0_bits_taskID(ReadController_io_ReadIn_0_bits_taskID),
    .io_ReadIn_1_ready(ReadController_io_ReadIn_1_ready),
    .io_ReadIn_1_valid(ReadController_io_ReadIn_1_valid),
    .io_ReadIn_1_bits_address(ReadController_io_ReadIn_1_bits_address),
    .io_ReadIn_1_bits_taskID(ReadController_io_ReadIn_1_bits_taskID),
    .io_ReadIn_2_ready(ReadController_io_ReadIn_2_ready),
    .io_ReadIn_2_valid(ReadController_io_ReadIn_2_valid),
    .io_ReadIn_2_bits_address(ReadController_io_ReadIn_2_bits_address),
    .io_ReadIn_2_bits_taskID(ReadController_io_ReadIn_2_bits_taskID),
    .io_ReadIn_3_ready(ReadController_io_ReadIn_3_ready),
    .io_ReadIn_3_valid(ReadController_io_ReadIn_3_valid),
    .io_ReadIn_3_bits_address(ReadController_io_ReadIn_3_bits_address),
    .io_ReadIn_3_bits_taskID(ReadController_io_ReadIn_3_bits_taskID),
    .io_ReadIn_4_ready(ReadController_io_ReadIn_4_ready),
    .io_ReadIn_4_valid(ReadController_io_ReadIn_4_valid),
    .io_ReadIn_4_bits_address(ReadController_io_ReadIn_4_bits_address),
    .io_ReadIn_4_bits_taskID(ReadController_io_ReadIn_4_bits_taskID),
    .io_ReadIn_5_ready(ReadController_io_ReadIn_5_ready),
    .io_ReadIn_5_valid(ReadController_io_ReadIn_5_valid),
    .io_ReadIn_5_bits_address(ReadController_io_ReadIn_5_bits_address),
    .io_ReadIn_5_bits_taskID(ReadController_io_ReadIn_5_bits_taskID),
    .io_ReadIn_6_ready(ReadController_io_ReadIn_6_ready),
    .io_ReadIn_6_valid(ReadController_io_ReadIn_6_valid),
    .io_ReadIn_6_bits_address(ReadController_io_ReadIn_6_bits_address),
    .io_ReadIn_6_bits_taskID(ReadController_io_ReadIn_6_bits_taskID),
    .io_ReadIn_7_ready(ReadController_io_ReadIn_7_ready),
    .io_ReadIn_7_valid(ReadController_io_ReadIn_7_valid),
    .io_ReadIn_7_bits_address(ReadController_io_ReadIn_7_bits_address),
    .io_ReadIn_7_bits_taskID(ReadController_io_ReadIn_7_bits_taskID),
    .io_ReadIn_8_ready(ReadController_io_ReadIn_8_ready),
    .io_ReadIn_8_valid(ReadController_io_ReadIn_8_valid),
    .io_ReadIn_8_bits_address(ReadController_io_ReadIn_8_bits_address),
    .io_ReadIn_8_bits_taskID(ReadController_io_ReadIn_8_bits_taskID),
    .io_ReadIn_9_ready(ReadController_io_ReadIn_9_ready),
    .io_ReadIn_9_valid(ReadController_io_ReadIn_9_valid),
    .io_ReadIn_9_bits_address(ReadController_io_ReadIn_9_bits_address),
    .io_ReadIn_9_bits_taskID(ReadController_io_ReadIn_9_bits_taskID),
    .io_ReadIn_10_ready(ReadController_io_ReadIn_10_ready),
    .io_ReadIn_10_valid(ReadController_io_ReadIn_10_valid),
    .io_ReadIn_10_bits_address(ReadController_io_ReadIn_10_bits_address),
    .io_ReadIn_10_bits_taskID(ReadController_io_ReadIn_10_bits_taskID),
    .io_ReadIn_11_ready(ReadController_io_ReadIn_11_ready),
    .io_ReadIn_11_valid(ReadController_io_ReadIn_11_valid),
    .io_ReadIn_11_bits_address(ReadController_io_ReadIn_11_bits_address),
    .io_ReadIn_11_bits_taskID(ReadController_io_ReadIn_11_bits_taskID),
    .io_ReadIn_12_ready(ReadController_io_ReadIn_12_ready),
    .io_ReadIn_12_valid(ReadController_io_ReadIn_12_valid),
    .io_ReadIn_12_bits_address(ReadController_io_ReadIn_12_bits_address),
    .io_ReadIn_12_bits_taskID(ReadController_io_ReadIn_12_bits_taskID),
    .io_ReadIn_13_ready(ReadController_io_ReadIn_13_ready),
    .io_ReadIn_13_valid(ReadController_io_ReadIn_13_valid),
    .io_ReadIn_13_bits_address(ReadController_io_ReadIn_13_bits_address),
    .io_ReadIn_13_bits_taskID(ReadController_io_ReadIn_13_bits_taskID),
    .io_ReadIn_14_ready(ReadController_io_ReadIn_14_ready),
    .io_ReadIn_14_valid(ReadController_io_ReadIn_14_valid),
    .io_ReadIn_14_bits_address(ReadController_io_ReadIn_14_bits_address),
    .io_ReadIn_14_bits_taskID(ReadController_io_ReadIn_14_bits_taskID),
    .io_ReadIn_15_ready(ReadController_io_ReadIn_15_ready),
    .io_ReadIn_15_valid(ReadController_io_ReadIn_15_valid),
    .io_ReadIn_15_bits_address(ReadController_io_ReadIn_15_bits_address),
    .io_ReadIn_15_bits_taskID(ReadController_io_ReadIn_15_bits_taskID),
    .io_ReadIn_16_ready(ReadController_io_ReadIn_16_ready),
    .io_ReadIn_16_valid(ReadController_io_ReadIn_16_valid),
    .io_ReadIn_16_bits_address(ReadController_io_ReadIn_16_bits_address),
    .io_ReadIn_16_bits_taskID(ReadController_io_ReadIn_16_bits_taskID),
    .io_ReadIn_17_ready(ReadController_io_ReadIn_17_ready),
    .io_ReadIn_17_valid(ReadController_io_ReadIn_17_valid),
    .io_ReadIn_17_bits_address(ReadController_io_ReadIn_17_bits_address),
    .io_ReadIn_17_bits_taskID(ReadController_io_ReadIn_17_bits_taskID),
    .io_ReadIn_18_ready(ReadController_io_ReadIn_18_ready),
    .io_ReadIn_18_valid(ReadController_io_ReadIn_18_valid),
    .io_ReadIn_18_bits_address(ReadController_io_ReadIn_18_bits_address),
    .io_ReadIn_18_bits_taskID(ReadController_io_ReadIn_18_bits_taskID),
    .io_ReadOut_0_valid(ReadController_io_ReadOut_0_valid),
    .io_ReadOut_0_data(ReadController_io_ReadOut_0_data),
    .io_ReadOut_1_valid(ReadController_io_ReadOut_1_valid),
    .io_ReadOut_1_data(ReadController_io_ReadOut_1_data),
    .io_ReadOut_2_valid(ReadController_io_ReadOut_2_valid),
    .io_ReadOut_2_data(ReadController_io_ReadOut_2_data),
    .io_ReadOut_3_valid(ReadController_io_ReadOut_3_valid),
    .io_ReadOut_3_data(ReadController_io_ReadOut_3_data),
    .io_ReadOut_4_valid(ReadController_io_ReadOut_4_valid),
    .io_ReadOut_4_data(ReadController_io_ReadOut_4_data),
    .io_ReadOut_5_valid(ReadController_io_ReadOut_5_valid),
    .io_ReadOut_5_data(ReadController_io_ReadOut_5_data),
    .io_ReadOut_6_valid(ReadController_io_ReadOut_6_valid),
    .io_ReadOut_6_data(ReadController_io_ReadOut_6_data),
    .io_ReadOut_7_valid(ReadController_io_ReadOut_7_valid),
    .io_ReadOut_7_data(ReadController_io_ReadOut_7_data),
    .io_ReadOut_8_valid(ReadController_io_ReadOut_8_valid),
    .io_ReadOut_8_data(ReadController_io_ReadOut_8_data),
    .io_ReadOut_9_valid(ReadController_io_ReadOut_9_valid),
    .io_ReadOut_9_data(ReadController_io_ReadOut_9_data),
    .io_ReadOut_10_valid(ReadController_io_ReadOut_10_valid),
    .io_ReadOut_10_data(ReadController_io_ReadOut_10_data),
    .io_ReadOut_11_valid(ReadController_io_ReadOut_11_valid),
    .io_ReadOut_11_data(ReadController_io_ReadOut_11_data),
    .io_ReadOut_12_valid(ReadController_io_ReadOut_12_valid),
    .io_ReadOut_12_data(ReadController_io_ReadOut_12_data),
    .io_ReadOut_13_valid(ReadController_io_ReadOut_13_valid),
    .io_ReadOut_13_data(ReadController_io_ReadOut_13_data),
    .io_ReadOut_14_valid(ReadController_io_ReadOut_14_valid),
    .io_ReadOut_14_data(ReadController_io_ReadOut_14_data),
    .io_ReadOut_15_valid(ReadController_io_ReadOut_15_valid),
    .io_ReadOut_15_data(ReadController_io_ReadOut_15_data),
    .io_ReadOut_16_valid(ReadController_io_ReadOut_16_valid),
    .io_ReadOut_16_data(ReadController_io_ReadOut_16_data),
    .io_ReadOut_17_valid(ReadController_io_ReadOut_17_valid),
    .io_ReadOut_17_data(ReadController_io_ReadOut_17_data),
    .io_ReadOut_18_valid(ReadController_io_ReadOut_18_valid),
    .io_ReadOut_18_data(ReadController_io_ReadOut_18_data),
    .io_MemReq_ready(ReadController_io_MemReq_ready),
    .io_MemReq_valid(ReadController_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadController_io_MemReq_bits_addr),
    .io_MemReq_bits_data(ReadController_io_MemReq_bits_data),
    .io_MemReq_bits_mask(ReadController_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(ReadController_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadController_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadController_io_MemReq_bits_iswrite),
    .io_MemResp_valid(ReadController_io_MemResp_valid),
    .io_MemResp_bits_data(ReadController_io_MemResp_bits_data),
    .io_MemResp_bits_tag(ReadController_io_MemResp_bits_tag)
  );
  ReadWriteArbiter ReadWriteArbiter ( // @[UnifiedController.scala 55:32]
    .clock(ReadWriteArbiter_clock),
    .io_ReadMemReq_ready(ReadWriteArbiter_io_ReadMemReq_ready),
    .io_ReadMemReq_valid(ReadWriteArbiter_io_ReadMemReq_valid),
    .io_ReadMemReq_bits_addr(ReadWriteArbiter_io_ReadMemReq_bits_addr),
    .io_ReadMemReq_bits_data(ReadWriteArbiter_io_ReadMemReq_bits_data),
    .io_ReadMemReq_bits_mask(ReadWriteArbiter_io_ReadMemReq_bits_mask),
    .io_ReadMemReq_bits_tag(ReadWriteArbiter_io_ReadMemReq_bits_tag),
    .io_ReadMemReq_bits_taskID(ReadWriteArbiter_io_ReadMemReq_bits_taskID),
    .io_ReadMemReq_bits_iswrite(ReadWriteArbiter_io_ReadMemReq_bits_iswrite),
    .io_WriteMemReq_ready(ReadWriteArbiter_io_WriteMemReq_ready),
    .io_WriteMemReq_valid(ReadWriteArbiter_io_WriteMemReq_valid),
    .io_WriteMemReq_bits_addr(ReadWriteArbiter_io_WriteMemReq_bits_addr),
    .io_WriteMemReq_bits_data(ReadWriteArbiter_io_WriteMemReq_bits_data),
    .io_WriteMemReq_bits_mask(ReadWriteArbiter_io_WriteMemReq_bits_mask),
    .io_WriteMemReq_bits_tag(ReadWriteArbiter_io_WriteMemReq_bits_tag),
    .io_WriteMemReq_bits_taskID(ReadWriteArbiter_io_WriteMemReq_bits_taskID),
    .io_WriteMemReq_bits_iswrite(ReadWriteArbiter_io_WriteMemReq_bits_iswrite),
    .io_MemResp_valid(ReadWriteArbiter_io_MemResp_valid),
    .io_MemResp_bits_data(ReadWriteArbiter_io_MemResp_bits_data),
    .io_MemResp_bits_tag(ReadWriteArbiter_io_MemResp_bits_tag),
    .io_MemResp_bits_iswrite(ReadWriteArbiter_io_MemResp_bits_iswrite),
    .io_ReadMemResp_valid(ReadWriteArbiter_io_ReadMemResp_valid),
    .io_ReadMemResp_bits_data(ReadWriteArbiter_io_ReadMemResp_bits_data),
    .io_ReadMemResp_bits_tag(ReadWriteArbiter_io_ReadMemResp_bits_tag),
    .io_WriteMemResp_valid(ReadWriteArbiter_io_WriteMemResp_valid),
    .io_WriteMemResp_bits_data(ReadWriteArbiter_io_WriteMemResp_bits_data),
    .io_WriteMemResp_bits_tag(ReadWriteArbiter_io_WriteMemResp_bits_tag),
    .io_MemReq_ready(ReadWriteArbiter_io_MemReq_ready),
    .io_MemReq_valid(ReadWriteArbiter_io_MemReq_valid),
    .io_MemReq_bits_addr(ReadWriteArbiter_io_MemReq_bits_addr),
    .io_MemReq_bits_data(ReadWriteArbiter_io_MemReq_bits_data),
    .io_MemReq_bits_mask(ReadWriteArbiter_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(ReadWriteArbiter_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(ReadWriteArbiter_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(ReadWriteArbiter_io_MemReq_bits_iswrite)
  );
  assign _T = io_MemReq_ready & io_MemReq_valid; // @[Decoupled.scala 40:37]
  assign _T_1 = $unsigned(reset); // @[UnifiedController.scala 92:15]
  assign _T_2 = _T_1 == 1'h0; // @[UnifiedController.scala 92:15]
  assign io_WriteIn_0_ready = WriteController_io_WriteIn_0_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteIn_1_ready = WriteController_io_WriteIn_1_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteIn_2_ready = WriteController_io_WriteIn_2_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteIn_3_ready = WriteController_io_WriteIn_3_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteIn_4_ready = WriteController_io_WriteIn_4_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteIn_5_ready = WriteController_io_WriteIn_5_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteIn_6_ready = WriteController_io_WriteIn_6_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteIn_7_ready = WriteController_io_WriteIn_7_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteIn_8_ready = WriteController_io_WriteIn_8_ready; // @[UnifiedController.scala 63:35]
  assign io_WriteOut_0_valid = WriteController_io_WriteOut_0_valid; // @[UnifiedController.scala 64:20]
  assign io_WriteOut_1_valid = WriteController_io_WriteOut_1_valid; // @[UnifiedController.scala 64:20]
  assign io_WriteOut_2_valid = WriteController_io_WriteOut_2_valid; // @[UnifiedController.scala 64:20]
  assign io_WriteOut_3_valid = WriteController_io_WriteOut_3_valid; // @[UnifiedController.scala 64:20]
  assign io_WriteOut_4_valid = WriteController_io_WriteOut_4_valid; // @[UnifiedController.scala 64:20]
  assign io_WriteOut_5_valid = WriteController_io_WriteOut_5_valid; // @[UnifiedController.scala 64:20]
  assign io_WriteOut_6_valid = WriteController_io_WriteOut_6_valid; // @[UnifiedController.scala 64:20]
  assign io_WriteOut_7_valid = WriteController_io_WriteOut_7_valid; // @[UnifiedController.scala 64:20]
  assign io_WriteOut_8_valid = WriteController_io_WriteOut_8_valid; // @[UnifiedController.scala 64:20]
  assign io_ReadIn_0_ready = ReadController_io_ReadIn_0_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_1_ready = ReadController_io_ReadIn_1_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_2_ready = ReadController_io_ReadIn_2_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_3_ready = ReadController_io_ReadIn_3_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_4_ready = ReadController_io_ReadIn_4_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_5_ready = ReadController_io_ReadIn_5_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_6_ready = ReadController_io_ReadIn_6_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_7_ready = ReadController_io_ReadIn_7_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_8_ready = ReadController_io_ReadIn_8_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_9_ready = ReadController_io_ReadIn_9_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_10_ready = ReadController_io_ReadIn_10_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_11_ready = ReadController_io_ReadIn_11_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_12_ready = ReadController_io_ReadIn_12_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_13_ready = ReadController_io_ReadIn_13_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_14_ready = ReadController_io_ReadIn_14_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_15_ready = ReadController_io_ReadIn_15_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_16_ready = ReadController_io_ReadIn_16_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_17_ready = ReadController_io_ReadIn_17_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadIn_18_ready = ReadController_io_ReadIn_18_ready; // @[UnifiedController.scala 69:33]
  assign io_ReadOut_0_valid = ReadController_io_ReadOut_0_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_0_data = ReadController_io_ReadOut_0_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_1_valid = ReadController_io_ReadOut_1_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_1_data = ReadController_io_ReadOut_1_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_2_valid = ReadController_io_ReadOut_2_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_2_data = ReadController_io_ReadOut_2_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_3_valid = ReadController_io_ReadOut_3_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_3_data = ReadController_io_ReadOut_3_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_4_valid = ReadController_io_ReadOut_4_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_4_data = ReadController_io_ReadOut_4_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_5_valid = ReadController_io_ReadOut_5_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_5_data = ReadController_io_ReadOut_5_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_6_valid = ReadController_io_ReadOut_6_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_6_data = ReadController_io_ReadOut_6_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_7_valid = ReadController_io_ReadOut_7_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_7_data = ReadController_io_ReadOut_7_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_8_valid = ReadController_io_ReadOut_8_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_8_data = ReadController_io_ReadOut_8_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_9_valid = ReadController_io_ReadOut_9_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_9_data = ReadController_io_ReadOut_9_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_10_valid = ReadController_io_ReadOut_10_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_10_data = ReadController_io_ReadOut_10_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_11_valid = ReadController_io_ReadOut_11_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_11_data = ReadController_io_ReadOut_11_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_12_valid = ReadController_io_ReadOut_12_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_12_data = ReadController_io_ReadOut_12_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_13_valid = ReadController_io_ReadOut_13_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_13_data = ReadController_io_ReadOut_13_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_14_valid = ReadController_io_ReadOut_14_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_14_data = ReadController_io_ReadOut_14_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_15_valid = ReadController_io_ReadOut_15_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_15_data = ReadController_io_ReadOut_15_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_16_valid = ReadController_io_ReadOut_16_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_16_data = ReadController_io_ReadOut_16_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_17_valid = ReadController_io_ReadOut_17_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_17_data = ReadController_io_ReadOut_17_data; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_18_valid = ReadController_io_ReadOut_18_valid; // @[UnifiedController.scala 70:19]
  assign io_ReadOut_18_data = ReadController_io_ReadOut_18_data; // @[UnifiedController.scala 70:19]
  assign io_MemReq_valid = ReadWriteArbiter_io_MemReq_valid; // @[UnifiedController.scala 83:19]
  assign io_MemReq_bits_addr = ReadWriteArbiter_io_MemReq_bits_addr; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_data = ReadWriteArbiter_io_MemReq_bits_data; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_mask = ReadWriteArbiter_io_MemReq_bits_mask; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_tag = ReadWriteArbiter_io_MemReq_bits_tag; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_taskID = ReadWriteArbiter_io_MemReq_bits_taskID; // @[UnifiedController.scala 82:18]
  assign io_MemReq_bits_iswrite = ReadWriteArbiter_io_MemReq_bits_iswrite; // @[UnifiedController.scala 82:18]
  assign WriteController_clock = clock;
  assign WriteController_reset = reset;
  assign WriteController_io_WriteIn_0_valid = io_WriteIn_0_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_0_bits_address = io_WriteIn_0_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_0_bits_data = io_WriteIn_0_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_0_bits_taskID = io_WriteIn_0_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_1_valid = io_WriteIn_1_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_1_bits_address = io_WriteIn_1_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_1_bits_data = io_WriteIn_1_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_1_bits_taskID = io_WriteIn_1_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_2_valid = io_WriteIn_2_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_2_bits_address = io_WriteIn_2_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_2_bits_data = io_WriteIn_2_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_2_bits_taskID = io_WriteIn_2_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_3_valid = io_WriteIn_3_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_3_bits_address = io_WriteIn_3_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_3_bits_data = io_WriteIn_3_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_3_bits_taskID = io_WriteIn_3_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_4_valid = io_WriteIn_4_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_4_bits_address = io_WriteIn_4_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_4_bits_data = io_WriteIn_4_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_4_bits_taskID = io_WriteIn_4_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_5_valid = io_WriteIn_5_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_5_bits_address = io_WriteIn_5_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_5_bits_data = io_WriteIn_5_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_5_bits_taskID = io_WriteIn_5_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_6_valid = io_WriteIn_6_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_6_bits_address = io_WriteIn_6_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_6_bits_data = io_WriteIn_6_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_6_bits_taskID = io_WriteIn_6_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_7_valid = io_WriteIn_7_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_7_bits_address = io_WriteIn_7_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_7_bits_data = io_WriteIn_7_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_7_bits_taskID = io_WriteIn_7_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_8_valid = io_WriteIn_8_valid; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_8_bits_address = io_WriteIn_8_bits_address; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_8_bits_data = io_WriteIn_8_bits_data; // @[UnifiedController.scala 63:35]
  assign WriteController_io_WriteIn_8_bits_taskID = io_WriteIn_8_bits_taskID; // @[UnifiedController.scala 63:35]
  assign WriteController_io_MemReq_ready = ReadWriteArbiter_io_WriteMemReq_ready; // @[UnifiedController.scala 77:35]
  assign WriteController_io_MemResp_valid = ReadWriteArbiter_io_WriteMemResp_valid; // @[UnifiedController.scala 78:30]
  assign WriteController_io_MemResp_bits_data = ReadWriteArbiter_io_WriteMemResp_bits_data; // @[UnifiedController.scala 78:30]
  assign WriteController_io_MemResp_bits_tag = ReadWriteArbiter_io_WriteMemResp_bits_tag; // @[UnifiedController.scala 78:30]
  assign ReadController_clock = clock;
  assign ReadController_reset = reset;
  assign ReadController_io_ReadIn_0_valid = io_ReadIn_0_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_0_bits_address = io_ReadIn_0_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_0_bits_taskID = io_ReadIn_0_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_1_valid = io_ReadIn_1_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_1_bits_address = io_ReadIn_1_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_1_bits_taskID = io_ReadIn_1_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_2_valid = io_ReadIn_2_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_2_bits_address = io_ReadIn_2_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_2_bits_taskID = io_ReadIn_2_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_3_valid = io_ReadIn_3_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_3_bits_address = io_ReadIn_3_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_3_bits_taskID = io_ReadIn_3_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_4_valid = io_ReadIn_4_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_4_bits_address = io_ReadIn_4_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_4_bits_taskID = io_ReadIn_4_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_5_valid = io_ReadIn_5_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_5_bits_address = io_ReadIn_5_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_5_bits_taskID = io_ReadIn_5_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_6_valid = io_ReadIn_6_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_6_bits_address = io_ReadIn_6_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_6_bits_taskID = io_ReadIn_6_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_7_valid = io_ReadIn_7_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_7_bits_address = io_ReadIn_7_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_7_bits_taskID = io_ReadIn_7_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_8_valid = io_ReadIn_8_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_8_bits_address = io_ReadIn_8_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_8_bits_taskID = io_ReadIn_8_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_9_valid = io_ReadIn_9_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_9_bits_address = io_ReadIn_9_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_9_bits_taskID = io_ReadIn_9_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_10_valid = io_ReadIn_10_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_10_bits_address = io_ReadIn_10_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_10_bits_taskID = io_ReadIn_10_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_11_valid = io_ReadIn_11_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_11_bits_address = io_ReadIn_11_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_11_bits_taskID = io_ReadIn_11_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_12_valid = io_ReadIn_12_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_12_bits_address = io_ReadIn_12_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_12_bits_taskID = io_ReadIn_12_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_13_valid = io_ReadIn_13_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_13_bits_address = io_ReadIn_13_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_13_bits_taskID = io_ReadIn_13_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_14_valid = io_ReadIn_14_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_14_bits_address = io_ReadIn_14_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_14_bits_taskID = io_ReadIn_14_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_15_valid = io_ReadIn_15_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_15_bits_address = io_ReadIn_15_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_15_bits_taskID = io_ReadIn_15_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_16_valid = io_ReadIn_16_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_16_bits_address = io_ReadIn_16_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_16_bits_taskID = io_ReadIn_16_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_17_valid = io_ReadIn_17_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_17_bits_address = io_ReadIn_17_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_17_bits_taskID = io_ReadIn_17_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_18_valid = io_ReadIn_18_valid; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_18_bits_address = io_ReadIn_18_bits_address; // @[UnifiedController.scala 69:33]
  assign ReadController_io_ReadIn_18_bits_taskID = io_ReadIn_18_bits_taskID; // @[UnifiedController.scala 69:33]
  assign ReadController_io_MemReq_ready = ReadWriteArbiter_io_ReadMemReq_ready; // @[UnifiedController.scala 74:34]
  assign ReadController_io_MemResp_valid = ReadWriteArbiter_io_ReadMemResp_valid; // @[UnifiedController.scala 75:29]
  assign ReadController_io_MemResp_bits_data = ReadWriteArbiter_io_ReadMemResp_bits_data; // @[UnifiedController.scala 75:29]
  assign ReadController_io_MemResp_bits_tag = ReadWriteArbiter_io_ReadMemResp_bits_tag; // @[UnifiedController.scala 75:29]
  assign ReadWriteArbiter_clock = clock;
  assign ReadWriteArbiter_io_ReadMemReq_valid = ReadController_io_MemReq_valid; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_addr = ReadController_io_MemReq_bits_addr; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_data = ReadController_io_MemReq_bits_data; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_mask = ReadController_io_MemReq_bits_mask; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_tag = ReadController_io_MemReq_bits_tag; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_taskID = ReadController_io_MemReq_bits_taskID; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_ReadMemReq_bits_iswrite = ReadController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 74:34]
  assign ReadWriteArbiter_io_WriteMemReq_valid = WriteController_io_MemReq_valid; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_addr = WriteController_io_MemReq_bits_addr; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_data = WriteController_io_MemReq_bits_data; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_mask = WriteController_io_MemReq_bits_mask; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_tag = WriteController_io_MemReq_bits_tag; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_taskID = WriteController_io_MemReq_bits_taskID; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_WriteMemReq_bits_iswrite = WriteController_io_MemReq_bits_iswrite; // @[UnifiedController.scala 77:35]
  assign ReadWriteArbiter_io_MemResp_valid = io_MemResp_valid; // @[UnifiedController.scala 84:31]
  assign ReadWriteArbiter_io_MemResp_bits_data = io_MemResp_bits_data; // @[UnifiedController.scala 84:31]
  assign ReadWriteArbiter_io_MemResp_bits_tag = io_MemResp_bits_tag; // @[UnifiedController.scala 84:31]
  assign ReadWriteArbiter_io_MemResp_bits_iswrite = io_MemResp_bits_iswrite; // @[UnifiedController.scala 84:31]
  assign ReadWriteArbiter_io_MemReq_ready = io_MemReq_ready; // @[UnifiedController.scala 81:36]
  assign _GEN_0 = _T & io_MemReq_bits_iswrite; // @[UnifiedController.scala 92:15]
  assign _GEN_1 = io_MemReq_bits_iswrite == 1'h0; // @[UnifiedController.scala 94:15]
  assign _GEN_2 = _T & _GEN_1; // @[UnifiedController.scala 94:15]
  assign _GEN_3 = io_MemResp_valid & io_MemResp_bits_iswrite; // @[UnifiedController.scala 100:15]
  assign _GEN_4 = io_MemResp_bits_iswrite == 1'h0; // @[UnifiedController.scala 102:15]
  assign _GEN_5 = io_MemResp_valid & _GEN_4; // @[UnifiedController.scala 102:15]
  always @(posedge clock) begin
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_0 & _T_2) begin
          $fwrite(32'h80000002,"[LOG] [MemController] [MemReq]: Addr: %d, Data: %d, IsWrite: ST\n",io_MemReq_bits_addr,io_MemReq_bits_data); // @[UnifiedController.scala 92:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_2 & _T_2) begin
          $fwrite(32'h80000002,"[LOG] [MemController] [MemReq]: Addr: %d, Data: %d, IsWrite: LD\n",io_MemReq_bits_addr,io_MemReq_bits_data); // @[UnifiedController.scala 94:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_3 & _T_2) begin
          $fwrite(32'h80000002,"[LOG] [MemController] [MemResp]: Data: %d, IsWrite: ST\n",io_MemResp_bits_data); // @[UnifiedController.scala 100:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_5 & _T_2) begin
          $fwrite(32'h80000002,"[LOG] [MemController] [MemResp]: Data: %d, IsWrite: LD\n",io_MemReq_bits_data); // @[UnifiedController.scala 102:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SplitCallNew(
  input         clock,
  input         reset,
  output        io_In_ready,
  input         io_In_valid,
  input  [4:0]  io_In_bits_enable_taskID,
  input         io_In_bits_enable_control,
  input  [31:0] io_In_bits_data_field5_data,
  input  [31:0] io_In_bits_data_field4_data,
  input  [31:0] io_In_bits_data_field3_data,
  input  [4:0]  io_In_bits_data_field2_taskID,
  input  [31:0] io_In_bits_data_field2_data,
  input         io_In_bits_data_field1_predicate,
  input  [4:0]  io_In_bits_data_field1_taskID,
  input  [31:0] io_In_bits_data_field1_data,
  input  [4:0]  io_In_bits_data_field0_taskID,
  input  [31:0] io_In_bits_data_field0_data,
  input         io_Out_enable_ready,
  output        io_Out_enable_valid,
  output [4:0]  io_Out_enable_bits_taskID,
  output        io_Out_enable_bits_control,
  input         io_Out_data_field5_0_ready,
  output        io_Out_data_field5_0_valid,
  output [31:0] io_Out_data_field5_0_bits_data,
  input         io_Out_data_field5_1_ready,
  output        io_Out_data_field5_1_valid,
  output [31:0] io_Out_data_field5_1_bits_data,
  input         io_Out_data_field4_0_ready,
  output        io_Out_data_field4_0_valid,
  output [31:0] io_Out_data_field4_0_bits_data,
  input         io_Out_data_field3_0_ready,
  output        io_Out_data_field3_0_valid,
  output [31:0] io_Out_data_field3_0_bits_data,
  input         io_Out_data_field2_0_ready,
  output        io_Out_data_field2_0_valid,
  output [4:0]  io_Out_data_field2_0_bits_taskID,
  output [31:0] io_Out_data_field2_0_bits_data,
  input         io_Out_data_field1_0_ready,
  output        io_Out_data_field1_0_valid,
  output        io_Out_data_field1_0_bits_predicate,
  output [4:0]  io_Out_data_field1_0_bits_taskID,
  output [31:0] io_Out_data_field1_0_bits_data,
  input         io_Out_data_field1_1_ready,
  output        io_Out_data_field1_1_valid,
  output [4:0]  io_Out_data_field1_1_bits_taskID,
  output [31:0] io_Out_data_field1_1_bits_data,
  input         io_Out_data_field1_2_ready,
  output        io_Out_data_field1_2_valid,
  output [4:0]  io_Out_data_field1_2_bits_taskID,
  output [31:0] io_Out_data_field1_2_bits_data,
  input         io_Out_data_field1_3_ready,
  output        io_Out_data_field1_3_valid,
  output [4:0]  io_Out_data_field1_3_bits_taskID,
  output [31:0] io_Out_data_field1_3_bits_data,
  input         io_Out_data_field1_4_ready,
  output        io_Out_data_field1_4_valid,
  output [4:0]  io_Out_data_field1_4_bits_taskID,
  output [31:0] io_Out_data_field1_4_bits_data,
  input         io_Out_data_field1_5_ready,
  output        io_Out_data_field1_5_valid,
  output [4:0]  io_Out_data_field1_5_bits_taskID,
  output [31:0] io_Out_data_field1_5_bits_data,
  input         io_Out_data_field1_6_ready,
  output        io_Out_data_field1_6_valid,
  output [4:0]  io_Out_data_field1_6_bits_taskID,
  output [31:0] io_Out_data_field1_6_bits_data,
  input         io_Out_data_field1_7_ready,
  output        io_Out_data_field1_7_valid,
  output [4:0]  io_Out_data_field1_7_bits_taskID,
  output [31:0] io_Out_data_field1_7_bits_data,
  input         io_Out_data_field1_8_ready,
  output        io_Out_data_field1_8_valid,
  output [4:0]  io_Out_data_field1_8_bits_taskID,
  output [31:0] io_Out_data_field1_8_bits_data,
  input         io_Out_data_field0_0_ready,
  output        io_Out_data_field0_0_valid,
  output [4:0]  io_Out_data_field0_0_bits_taskID,
  output [31:0] io_Out_data_field0_0_bits_data
);
  reg [4:0] inputReg_enable_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_0;
  reg  inputReg_enable_control; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_1;
  reg [31:0] inputReg_data_field5_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_2;
  reg [31:0] inputReg_data_field4_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_3;
  reg [31:0] inputReg_data_field3_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_4;
  reg [4:0] inputReg_data_field2_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_5;
  reg [31:0] inputReg_data_field2_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_6;
  reg  inputReg_data_field1_predicate; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_7;
  reg [4:0] inputReg_data_field1_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_8;
  reg [31:0] inputReg_data_field1_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_9;
  reg [4:0] inputReg_data_field0_taskID; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_10;
  reg [31:0] inputReg_data_field0_data; // @[SplitDecoupled.scala 152:26]
  reg [31:0] _RAND_11;
  reg  enableValidReg; // @[SplitDecoupled.scala 154:31]
  reg [31:0] _RAND_12;
  reg  allValid_0; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_13;
  reg  outputValidReg_1_0; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_14;
  reg  outputValidReg_1_1; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_15;
  reg  outputValidReg_1_2; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_16;
  reg  outputValidReg_1_3; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_17;
  reg  outputValidReg_1_4; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_18;
  reg  outputValidReg_1_5; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_19;
  reg  outputValidReg_1_6; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_20;
  reg  outputValidReg_1_7; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_21;
  reg  outputValidReg_1_8; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_22;
  reg  allValid_2; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_23;
  reg  allValid_3; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_24;
  reg  allValid_4; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_25;
  reg  outputValidReg_5_0; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_26;
  reg  outputValidReg_5_1; // @[SplitDecoupled.scala 157:49]
  reg [31:0] _RAND_27;
  wire  _T_22; // @[SplitDecoupled.scala 161:51]
  wire  _T_23; // @[SplitDecoupled.scala 161:51]
  wire  _T_24; // @[SplitDecoupled.scala 161:51]
  wire  _T_25; // @[SplitDecoupled.scala 161:51]
  wire  _T_26; // @[SplitDecoupled.scala 161:51]
  wire  _T_27; // @[SplitDecoupled.scala 161:51]
  wire  _T_28; // @[SplitDecoupled.scala 161:51]
  wire  allValid_1; // @[SplitDecoupled.scala 161:51]
  wire  allValid_5; // @[SplitDecoupled.scala 161:51]
  reg  state; // @[SplitDecoupled.scala 166:22]
  reg [31:0] _RAND_28;
  wire  _T_29; // @[SplitDecoupled.scala 168:24]
  wire  _T_30; // @[Conditional.scala 37:30]
  wire  _T_31; // @[Decoupled.scala 40:37]
  wire  _GEN_0; // @[SplitDecoupled.scala 172:27]
  wire  _T_33; // @[SplitDecoupled.scala 178:36]
  wire  _T_34; // @[SplitDecoupled.scala 178:36]
  wire  _T_35; // @[SplitDecoupled.scala 178:36]
  wire  _T_36; // @[SplitDecoupled.scala 178:36]
  wire  _T_37; // @[SplitDecoupled.scala 178:36]
  wire  _T_38; // @[SplitDecoupled.scala 178:13]
  wire  _T_39; // @[SplitDecoupled.scala 178:45]
  wire  _T_40; // @[SplitDecoupled.scala 178:42]
  wire  _T_42; // @[SplitDecoupled.scala 186:24]
  wire  _GEN_44; // @[SplitDecoupled.scala 186:45]
  wire  _T_44; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_46; // @[SplitDecoupled.scala 186:45]
  wire  _T_48; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_48; // @[SplitDecoupled.scala 186:45]
  wire  _T_52; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_50; // @[SplitDecoupled.scala 186:45]
  wire  _T_56; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_52; // @[SplitDecoupled.scala 186:45]
  wire  _T_60; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_54; // @[SplitDecoupled.scala 186:45]
  wire  _T_64; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_56; // @[SplitDecoupled.scala 186:45]
  wire  _T_68; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_58; // @[SplitDecoupled.scala 186:45]
  wire  _T_72; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_60; // @[SplitDecoupled.scala 186:45]
  wire  _T_76; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_62; // @[SplitDecoupled.scala 186:45]
  wire  _T_80; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_64; // @[SplitDecoupled.scala 186:45]
  wire  _T_84; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_66; // @[SplitDecoupled.scala 186:45]
  wire  _T_88; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_68; // @[SplitDecoupled.scala 186:45]
  wire  _T_92; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_70; // @[SplitDecoupled.scala 186:45]
  wire  _T_96; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_72; // @[SplitDecoupled.scala 186:45]
  wire  _T_100; // @[SplitDecoupled.scala 189:32]
  wire  _GEN_74; // @[SplitDecoupled.scala 197:41]
  wire  _T_104; // @[SplitDecoupled.scala 200:28]
  assign _T_22 = outputValidReg_1_0 | outputValidReg_1_1; // @[SplitDecoupled.scala 161:51]
  assign _T_23 = _T_22 | outputValidReg_1_2; // @[SplitDecoupled.scala 161:51]
  assign _T_24 = _T_23 | outputValidReg_1_3; // @[SplitDecoupled.scala 161:51]
  assign _T_25 = _T_24 | outputValidReg_1_4; // @[SplitDecoupled.scala 161:51]
  assign _T_26 = _T_25 | outputValidReg_1_5; // @[SplitDecoupled.scala 161:51]
  assign _T_27 = _T_26 | outputValidReg_1_6; // @[SplitDecoupled.scala 161:51]
  assign _T_28 = _T_27 | outputValidReg_1_7; // @[SplitDecoupled.scala 161:51]
  assign allValid_1 = _T_28 | outputValidReg_1_8; // @[SplitDecoupled.scala 161:51]
  assign allValid_5 = outputValidReg_5_0 | outputValidReg_5_1; // @[SplitDecoupled.scala 161:51]
  assign _T_29 = state == 1'h0; // @[SplitDecoupled.scala 168:24]
  assign _T_30 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_31 = io_In_ready & io_In_valid; // @[Decoupled.scala 40:37]
  assign _GEN_0 = _T_31 | state; // @[SplitDecoupled.scala 172:27]
  assign _T_33 = allValid_0 | allValid_1; // @[SplitDecoupled.scala 178:36]
  assign _T_34 = _T_33 | allValid_2; // @[SplitDecoupled.scala 178:36]
  assign _T_35 = _T_34 | allValid_3; // @[SplitDecoupled.scala 178:36]
  assign _T_36 = _T_35 | allValid_4; // @[SplitDecoupled.scala 178:36]
  assign _T_37 = _T_36 | allValid_5; // @[SplitDecoupled.scala 178:36]
  assign _T_38 = _T_37 == 1'h0; // @[SplitDecoupled.scala 178:13]
  assign _T_39 = enableValidReg == 1'h0; // @[SplitDecoupled.scala 178:45]
  assign _T_40 = _T_38 & _T_39; // @[SplitDecoupled.scala 178:42]
  assign _T_42 = io_In_valid & _T_29; // @[SplitDecoupled.scala 186:24]
  assign _GEN_44 = _T_42 | allValid_0; // @[SplitDecoupled.scala 186:45]
  assign _T_44 = state & io_Out_data_field0_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_46 = _T_42 | outputValidReg_1_0; // @[SplitDecoupled.scala 186:45]
  assign _T_48 = state & io_Out_data_field1_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_48 = _T_42 | outputValidReg_1_1; // @[SplitDecoupled.scala 186:45]
  assign _T_52 = state & io_Out_data_field1_1_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_50 = _T_42 | outputValidReg_1_2; // @[SplitDecoupled.scala 186:45]
  assign _T_56 = state & io_Out_data_field1_2_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_52 = _T_42 | outputValidReg_1_3; // @[SplitDecoupled.scala 186:45]
  assign _T_60 = state & io_Out_data_field1_3_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_54 = _T_42 | outputValidReg_1_4; // @[SplitDecoupled.scala 186:45]
  assign _T_64 = state & io_Out_data_field1_4_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_56 = _T_42 | outputValidReg_1_5; // @[SplitDecoupled.scala 186:45]
  assign _T_68 = state & io_Out_data_field1_5_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_58 = _T_42 | outputValidReg_1_6; // @[SplitDecoupled.scala 186:45]
  assign _T_72 = state & io_Out_data_field1_6_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_60 = _T_42 | outputValidReg_1_7; // @[SplitDecoupled.scala 186:45]
  assign _T_76 = state & io_Out_data_field1_7_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_62 = _T_42 | outputValidReg_1_8; // @[SplitDecoupled.scala 186:45]
  assign _T_80 = state & io_Out_data_field1_8_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_64 = _T_42 | allValid_2; // @[SplitDecoupled.scala 186:45]
  assign _T_84 = state & io_Out_data_field2_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_66 = _T_42 | allValid_3; // @[SplitDecoupled.scala 186:45]
  assign _T_88 = state & io_Out_data_field3_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_68 = _T_42 | allValid_4; // @[SplitDecoupled.scala 186:45]
  assign _T_92 = state & io_Out_data_field4_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_70 = _T_42 | outputValidReg_5_0; // @[SplitDecoupled.scala 186:45]
  assign _T_96 = state & io_Out_data_field5_0_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_72 = _T_42 | outputValidReg_5_1; // @[SplitDecoupled.scala 186:45]
  assign _T_100 = state & io_Out_data_field5_1_ready; // @[SplitDecoupled.scala 189:32]
  assign _GEN_74 = _T_42 | enableValidReg; // @[SplitDecoupled.scala 197:41]
  assign _T_104 = state & io_Out_enable_ready; // @[SplitDecoupled.scala 200:28]
  assign io_In_ready = state == 1'h0; // @[SplitDecoupled.scala 168:15]
  assign io_Out_enable_valid = enableValidReg; // @[SplitDecoupled.scala 203:23]
  assign io_Out_enable_bits_taskID = inputReg_enable_taskID; // @[SplitDecoupled.scala 204:22]
  assign io_Out_enable_bits_control = inputReg_enable_control; // @[SplitDecoupled.scala 204:22]
  assign io_Out_data_field5_0_valid = outputValidReg_5_0; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field5_0_bits_data = inputReg_data_field5_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field5_1_valid = outputValidReg_5_1; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field5_1_bits_data = inputReg_data_field5_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field4_0_valid = allValid_4; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field4_0_bits_data = inputReg_data_field4_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field3_0_valid = allValid_3; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field3_0_bits_data = inputReg_data_field3_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field2_0_valid = allValid_2; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field2_0_bits_taskID = inputReg_data_field2_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field2_0_bits_data = inputReg_data_field2_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_0_valid = outputValidReg_1_0; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_0_bits_predicate = inputReg_data_field1_predicate; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_0_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_0_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_1_valid = outputValidReg_1_1; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_1_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_1_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_2_valid = outputValidReg_1_2; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_2_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_2_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_3_valid = outputValidReg_1_3; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_3_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_3_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_4_valid = outputValidReg_1_4; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_4_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_4_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_5_valid = outputValidReg_1_5; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_5_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_5_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_6_valid = outputValidReg_1_6; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_6_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_6_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_7_valid = outputValidReg_1_7; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_7_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_7_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_8_valid = outputValidReg_1_8; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field1_8_bits_taskID = inputReg_data_field1_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field1_8_bits_data = inputReg_data_field1_data; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field0_0_valid = allValid_0; // @[SplitDecoupled.scala 192:40]
  assign io_Out_data_field0_0_bits_taskID = inputReg_data_field0_taskID; // @[SplitDecoupled.scala 193:39]
  assign io_Out_data_field0_0_bits_data = inputReg_data_field0_data; // @[SplitDecoupled.scala 193:39]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inputReg_enable_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inputReg_enable_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inputReg_data_field5_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  inputReg_data_field4_data = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  inputReg_data_field3_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  inputReg_data_field2_taskID = _RAND_5[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  inputReg_data_field2_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  inputReg_data_field1_predicate = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  inputReg_data_field1_taskID = _RAND_8[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  inputReg_data_field1_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  inputReg_data_field0_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  inputReg_data_field0_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  enableValidReg = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  allValid_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  outputValidReg_1_0 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  outputValidReg_1_1 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  outputValidReg_1_2 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  outputValidReg_1_3 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  outputValidReg_1_4 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  outputValidReg_1_5 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  outputValidReg_1_6 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  outputValidReg_1_7 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  outputValidReg_1_8 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  allValid_2 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  allValid_3 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  allValid_4 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  outputValidReg_5_0 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  outputValidReg_5_1 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  state = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      inputReg_enable_taskID <= 5'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_enable_taskID <= io_In_bits_enable_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_enable_control <= 1'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_enable_control <= io_In_bits_enable_control;
        end
      end
    end
    if (reset) begin
      inputReg_data_field5_data <= 32'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field5_data <= io_In_bits_data_field5_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field4_data <= 32'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field4_data <= io_In_bits_data_field4_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field3_data <= 32'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field3_data <= io_In_bits_data_field3_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field2_taskID <= 5'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field2_taskID <= io_In_bits_data_field2_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field2_data <= 32'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field2_data <= io_In_bits_data_field2_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field1_predicate <= 1'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field1_predicate <= io_In_bits_data_field1_predicate;
        end
      end
    end
    if (reset) begin
      inputReg_data_field1_taskID <= 5'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field1_taskID <= io_In_bits_data_field1_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field1_data <= 32'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field1_data <= io_In_bits_data_field1_data;
        end
      end
    end
    if (reset) begin
      inputReg_data_field0_taskID <= 5'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field0_taskID <= io_In_bits_data_field0_taskID;
        end
      end
    end
    if (reset) begin
      inputReg_data_field0_data <= 32'h0;
    end else begin
      if (_T_30) begin
        if (_T_31) begin
          inputReg_data_field0_data <= io_In_bits_data_field0_data;
        end
      end
    end
    if (reset) begin
      enableValidReg <= 1'h0;
    end else begin
      if (_T_104) begin
        enableValidReg <= 1'h0;
      end else begin
        enableValidReg <= _GEN_74;
      end
    end
    if (reset) begin
      allValid_0 <= 1'h0;
    end else begin
      if (_T_44) begin
        allValid_0 <= 1'h0;
      end else begin
        allValid_0 <= _GEN_44;
      end
    end
    if (reset) begin
      outputValidReg_1_0 <= 1'h0;
    end else begin
      if (_T_48) begin
        outputValidReg_1_0 <= 1'h0;
      end else begin
        outputValidReg_1_0 <= _GEN_46;
      end
    end
    if (reset) begin
      outputValidReg_1_1 <= 1'h0;
    end else begin
      if (_T_52) begin
        outputValidReg_1_1 <= 1'h0;
      end else begin
        outputValidReg_1_1 <= _GEN_48;
      end
    end
    if (reset) begin
      outputValidReg_1_2 <= 1'h0;
    end else begin
      if (_T_56) begin
        outputValidReg_1_2 <= 1'h0;
      end else begin
        outputValidReg_1_2 <= _GEN_50;
      end
    end
    if (reset) begin
      outputValidReg_1_3 <= 1'h0;
    end else begin
      if (_T_60) begin
        outputValidReg_1_3 <= 1'h0;
      end else begin
        outputValidReg_1_3 <= _GEN_52;
      end
    end
    if (reset) begin
      outputValidReg_1_4 <= 1'h0;
    end else begin
      if (_T_64) begin
        outputValidReg_1_4 <= 1'h0;
      end else begin
        outputValidReg_1_4 <= _GEN_54;
      end
    end
    if (reset) begin
      outputValidReg_1_5 <= 1'h0;
    end else begin
      if (_T_68) begin
        outputValidReg_1_5 <= 1'h0;
      end else begin
        outputValidReg_1_5 <= _GEN_56;
      end
    end
    if (reset) begin
      outputValidReg_1_6 <= 1'h0;
    end else begin
      if (_T_72) begin
        outputValidReg_1_6 <= 1'h0;
      end else begin
        outputValidReg_1_6 <= _GEN_58;
      end
    end
    if (reset) begin
      outputValidReg_1_7 <= 1'h0;
    end else begin
      if (_T_76) begin
        outputValidReg_1_7 <= 1'h0;
      end else begin
        outputValidReg_1_7 <= _GEN_60;
      end
    end
    if (reset) begin
      outputValidReg_1_8 <= 1'h0;
    end else begin
      if (_T_80) begin
        outputValidReg_1_8 <= 1'h0;
      end else begin
        outputValidReg_1_8 <= _GEN_62;
      end
    end
    if (reset) begin
      allValid_2 <= 1'h0;
    end else begin
      if (_T_84) begin
        allValid_2 <= 1'h0;
      end else begin
        allValid_2 <= _GEN_64;
      end
    end
    if (reset) begin
      allValid_3 <= 1'h0;
    end else begin
      if (_T_88) begin
        allValid_3 <= 1'h0;
      end else begin
        allValid_3 <= _GEN_66;
      end
    end
    if (reset) begin
      allValid_4 <= 1'h0;
    end else begin
      if (_T_92) begin
        allValid_4 <= 1'h0;
      end else begin
        allValid_4 <= _GEN_68;
      end
    end
    if (reset) begin
      outputValidReg_5_0 <= 1'h0;
    end else begin
      if (_T_96) begin
        outputValidReg_5_0 <= 1'h0;
      end else begin
        outputValidReg_5_0 <= _GEN_70;
      end
    end
    if (reset) begin
      outputValidReg_5_1 <= 1'h0;
    end else begin
      if (_T_100) begin
        outputValidReg_5_1 <= 1'h0;
      end else begin
        outputValidReg_5_1 <= _GEN_72;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_30) begin
        state <= _GEN_0;
      end else begin
        if (state) begin
          if (_T_40) begin
            state <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module LoopBlockNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input  [31:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input         io_InLiveIn_4_bits_predicate,
  input  [4:0]  io_InLiveIn_4_bits_taskID,
  input  [31:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input  [31:0] io_InLiveIn_5_bits_data,
  output        io_InLiveIn_6_ready,
  input         io_InLiveIn_6_valid,
  input         io_InLiveIn_6_bits_predicate,
  input  [4:0]  io_InLiveIn_6_bits_taskID,
  input  [31:0] io_InLiveIn_6_bits_data,
  output        io_InLiveIn_7_ready,
  input         io_InLiveIn_7_valid,
  input         io_InLiveIn_7_bits_predicate,
  input  [4:0]  io_InLiveIn_7_bits_taskID,
  input  [31:0] io_InLiveIn_7_bits_data,
  output        io_InLiveIn_8_ready,
  input         io_InLiveIn_8_valid,
  input         io_InLiveIn_8_bits_predicate,
  input  [4:0]  io_InLiveIn_8_bits_taskID,
  input  [31:0] io_InLiveIn_8_bits_data,
  output        io_InLiveIn_9_ready,
  input         io_InLiveIn_9_valid,
  input         io_InLiveIn_9_bits_predicate,
  input  [4:0]  io_InLiveIn_9_bits_taskID,
  input  [31:0] io_InLiveIn_9_bits_data,
  output        io_InLiveIn_10_ready,
  input         io_InLiveIn_10_valid,
  input  [4:0]  io_InLiveIn_10_bits_taskID,
  input  [31:0] io_InLiveIn_10_bits_data,
  output        io_InLiveIn_11_ready,
  input         io_InLiveIn_11_valid,
  input  [4:0]  io_InLiveIn_11_bits_taskID,
  input  [31:0] io_InLiveIn_11_bits_data,
  output        io_InLiveIn_12_ready,
  input         io_InLiveIn_12_valid,
  input         io_InLiveIn_12_bits_predicate,
  input  [4:0]  io_InLiveIn_12_bits_taskID,
  input  [31:0] io_InLiveIn_12_bits_data,
  output        io_InLiveIn_13_ready,
  input         io_InLiveIn_13_valid,
  input         io_InLiveIn_13_bits_predicate,
  input  [4:0]  io_InLiveIn_13_bits_taskID,
  input  [31:0] io_InLiveIn_13_bits_data,
  output        io_InLiveIn_14_ready,
  input         io_InLiveIn_14_valid,
  input         io_InLiveIn_14_bits_predicate,
  input  [4:0]  io_InLiveIn_14_bits_taskID,
  input  [31:0] io_InLiveIn_14_bits_data,
  output        io_InLiveIn_15_ready,
  input         io_InLiveIn_15_valid,
  input         io_InLiveIn_15_bits_predicate,
  input  [4:0]  io_InLiveIn_15_bits_taskID,
  input  [31:0] io_InLiveIn_15_bits_data,
  input         io_OutLiveIn_field15_0_ready,
  output        io_OutLiveIn_field15_0_valid,
  output        io_OutLiveIn_field15_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field15_0_bits_taskID,
  output [31:0] io_OutLiveIn_field15_0_bits_data,
  input         io_OutLiveIn_field14_0_ready,
  output        io_OutLiveIn_field14_0_valid,
  output        io_OutLiveIn_field14_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field14_0_bits_taskID,
  output [31:0] io_OutLiveIn_field14_0_bits_data,
  input         io_OutLiveIn_field13_0_ready,
  output        io_OutLiveIn_field13_0_valid,
  output        io_OutLiveIn_field13_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field13_0_bits_taskID,
  output [31:0] io_OutLiveIn_field13_0_bits_data,
  input         io_OutLiveIn_field12_0_ready,
  output        io_OutLiveIn_field12_0_valid,
  output        io_OutLiveIn_field12_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field12_0_bits_taskID,
  output [31:0] io_OutLiveIn_field12_0_bits_data,
  input         io_OutLiveIn_field11_0_ready,
  output        io_OutLiveIn_field11_0_valid,
  output [4:0]  io_OutLiveIn_field11_0_bits_taskID,
  output [31:0] io_OutLiveIn_field11_0_bits_data,
  input         io_OutLiveIn_field10_0_ready,
  output        io_OutLiveIn_field10_0_valid,
  output [4:0]  io_OutLiveIn_field10_0_bits_taskID,
  output [31:0] io_OutLiveIn_field10_0_bits_data,
  input         io_OutLiveIn_field10_1_ready,
  output        io_OutLiveIn_field10_1_valid,
  output [4:0]  io_OutLiveIn_field10_1_bits_taskID,
  output [31:0] io_OutLiveIn_field10_1_bits_data,
  input         io_OutLiveIn_field10_2_ready,
  output        io_OutLiveIn_field10_2_valid,
  output [4:0]  io_OutLiveIn_field10_2_bits_taskID,
  output [31:0] io_OutLiveIn_field10_2_bits_data,
  input         io_OutLiveIn_field10_3_ready,
  output        io_OutLiveIn_field10_3_valid,
  output [4:0]  io_OutLiveIn_field10_3_bits_taskID,
  output [31:0] io_OutLiveIn_field10_3_bits_data,
  input         io_OutLiveIn_field10_4_ready,
  output        io_OutLiveIn_field10_4_valid,
  output [4:0]  io_OutLiveIn_field10_4_bits_taskID,
  output [31:0] io_OutLiveIn_field10_4_bits_data,
  input         io_OutLiveIn_field10_5_ready,
  output        io_OutLiveIn_field10_5_valid,
  output [4:0]  io_OutLiveIn_field10_5_bits_taskID,
  output [31:0] io_OutLiveIn_field10_5_bits_data,
  input         io_OutLiveIn_field10_6_ready,
  output        io_OutLiveIn_field10_6_valid,
  output [4:0]  io_OutLiveIn_field10_6_bits_taskID,
  output [31:0] io_OutLiveIn_field10_6_bits_data,
  input         io_OutLiveIn_field10_7_ready,
  output        io_OutLiveIn_field10_7_valid,
  output [4:0]  io_OutLiveIn_field10_7_bits_taskID,
  output [31:0] io_OutLiveIn_field10_7_bits_data,
  input         io_OutLiveIn_field10_8_ready,
  output        io_OutLiveIn_field10_8_valid,
  output [4:0]  io_OutLiveIn_field10_8_bits_taskID,
  output [31:0] io_OutLiveIn_field10_8_bits_data,
  input         io_OutLiveIn_field9_0_ready,
  output        io_OutLiveIn_field9_0_valid,
  output        io_OutLiveIn_field9_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field9_0_bits_taskID,
  output [31:0] io_OutLiveIn_field9_0_bits_data,
  input         io_OutLiveIn_field8_0_ready,
  output        io_OutLiveIn_field8_0_valid,
  output        io_OutLiveIn_field8_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field8_0_bits_taskID,
  output [31:0] io_OutLiveIn_field8_0_bits_data,
  input         io_OutLiveIn_field7_0_ready,
  output        io_OutLiveIn_field7_0_valid,
  output        io_OutLiveIn_field7_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field7_0_bits_taskID,
  output [31:0] io_OutLiveIn_field7_0_bits_data,
  input         io_OutLiveIn_field6_0_ready,
  output        io_OutLiveIn_field6_0_valid,
  output        io_OutLiveIn_field6_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field6_0_bits_taskID,
  output [31:0] io_OutLiveIn_field6_0_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output [31:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output        io_OutLiveIn_field4_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field4_0_bits_taskID,
  output [31:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_2;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_3;
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_5;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_6;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_7;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_8;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg  in_live_in_R_4_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [4:0] in_live_in_R_4_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg [31:0] in_live_in_R_4_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_15;
  reg [31:0] in_live_in_R_5_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_16;
  reg  in_live_in_R_6_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_17;
  reg [4:0] in_live_in_R_6_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_18;
  reg [31:0] in_live_in_R_6_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_19;
  reg  in_live_in_R_7_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_20;
  reg [4:0] in_live_in_R_7_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_21;
  reg [31:0] in_live_in_R_7_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_22;
  reg  in_live_in_R_8_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_23;
  reg [4:0] in_live_in_R_8_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_24;
  reg [31:0] in_live_in_R_8_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_25;
  reg  in_live_in_R_9_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_26;
  reg [4:0] in_live_in_R_9_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_27;
  reg [31:0] in_live_in_R_9_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_28;
  reg [4:0] in_live_in_R_10_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_29;
  reg [31:0] in_live_in_R_10_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_30;
  reg [4:0] in_live_in_R_11_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_31;
  reg [31:0] in_live_in_R_11_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_32;
  reg  in_live_in_R_12_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_33;
  reg [4:0] in_live_in_R_12_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_34;
  reg [31:0] in_live_in_R_12_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_35;
  reg  in_live_in_R_13_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_36;
  reg [4:0] in_live_in_R_13_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_37;
  reg [31:0] in_live_in_R_13_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_38;
  reg  in_live_in_R_14_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_39;
  reg [4:0] in_live_in_R_14_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_40;
  reg [31:0] in_live_in_R_14_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_41;
  reg  in_live_in_R_15_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_42;
  reg [4:0] in_live_in_R_15_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_43;
  reg [31:0] in_live_in_R_15_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_44;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_45;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_46;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_47;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_48;
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_49;
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_50;
  reg  in_live_in_valid_R_6; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_51;
  reg  in_live_in_valid_R_7; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_52;
  reg  in_live_in_valid_R_8; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_53;
  reg  in_live_in_valid_R_9; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_54;
  reg  in_live_in_valid_R_10; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_55;
  reg  in_live_in_valid_R_11; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_56;
  reg  in_live_in_valid_R_12; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_57;
  reg  in_live_in_valid_R_13; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_58;
  reg  in_live_in_valid_R_14; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_59;
  reg  in_live_in_valid_R_15; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_60;
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_61;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_62;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_63;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_64;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_65;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_66;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_67;
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_68;
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_69;
  reg  out_live_in_valid_R_6_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_70;
  reg  out_live_in_valid_R_7_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_71;
  reg  out_live_in_valid_R_8_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_72;
  reg  out_live_in_valid_R_9_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_73;
  reg  out_live_in_valid_R_10_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_74;
  reg  out_live_in_valid_R_10_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_75;
  reg  out_live_in_valid_R_10_2; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_76;
  reg  out_live_in_valid_R_10_3; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_77;
  reg  out_live_in_valid_R_10_4; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_78;
  reg  out_live_in_valid_R_10_5; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_79;
  reg  out_live_in_valid_R_10_6; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_80;
  reg  out_live_in_valid_R_10_7; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_81;
  reg  out_live_in_valid_R_10_8; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_82;
  reg  out_live_in_valid_R_11_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_83;
  reg  out_live_in_valid_R_12_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_84;
  reg  out_live_in_valid_R_13_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_85;
  reg  out_live_in_valid_R_14_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_86;
  reg  out_live_in_valid_R_15_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_87;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_88;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_89;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_90;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_91;
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_92;
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_93;
  reg  out_live_in_fire_R_6_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_94;
  reg  out_live_in_fire_R_7_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_95;
  reg  out_live_in_fire_R_8_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_96;
  reg  out_live_in_fire_R_9_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_97;
  reg  out_live_in_fire_R_10_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_98;
  reg  out_live_in_fire_R_10_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_99;
  reg  out_live_in_fire_R_10_2; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_100;
  reg  out_live_in_fire_R_10_3; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_101;
  reg  out_live_in_fire_R_10_4; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_102;
  reg  out_live_in_fire_R_10_5; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_103;
  reg  out_live_in_fire_R_10_6; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_104;
  reg  out_live_in_fire_R_10_7; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_105;
  reg  out_live_in_fire_R_10_8; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_106;
  reg  out_live_in_fire_R_11_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_107;
  reg  out_live_in_fire_R_12_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_108;
  reg  out_live_in_fire_R_13_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_109;
  reg  out_live_in_fire_R_14_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_110;
  reg  out_live_in_fire_R_15_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_111;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_112;
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_113;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_114;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_115;
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_116;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_117;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_118;
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_119;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_120;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_121;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_122;
  wire  _T_28; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[LoopBlock.scala 603:33]
  wire [4:0] _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_32; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_34; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_36; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_38; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_40; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_42; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[LoopBlock.scala 623:33]
  wire  _T_44; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[LoopBlock.scala 623:33]
  wire  _T_46; // @[Decoupled.scala 40:37]
  wire  _GEN_37; // @[LoopBlock.scala 623:33]
  wire  _T_48; // @[Decoupled.scala 40:37]
  wire  _GEN_41; // @[LoopBlock.scala 623:33]
  wire  _T_50; // @[Decoupled.scala 40:37]
  wire  _GEN_45; // @[LoopBlock.scala 623:33]
  wire  _T_52; // @[Decoupled.scala 40:37]
  wire  _GEN_49; // @[LoopBlock.scala 623:33]
  wire  _T_54; // @[Decoupled.scala 40:37]
  wire  _GEN_53; // @[LoopBlock.scala 623:33]
  wire  _T_56; // @[Decoupled.scala 40:37]
  wire  _GEN_57; // @[LoopBlock.scala 623:33]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire  _GEN_61; // @[LoopBlock.scala 623:33]
  wire  _T_60; // @[Decoupled.scala 40:37]
  wire  _GEN_65; // @[LoopBlock.scala 623:33]
  wire  _T_62; // @[Decoupled.scala 40:37]
  wire  _GEN_69; // @[LoopBlock.scala 623:33]
  wire  _T_64; // @[Decoupled.scala 40:37]
  wire  _GEN_73; // @[LoopBlock.scala 623:33]
  wire  _T_66; // @[Decoupled.scala 40:37]
  wire  _GEN_77; // @[LoopBlock.scala 641:37]
  wire  _T_67; // @[Decoupled.scala 40:37]
  wire  _GEN_78; // @[LoopBlock.scala 704:39]
  wire  _T_68; // @[Decoupled.scala 40:37]
  wire  _GEN_79; // @[LoopBlock.scala 708:38]
  wire  _T_69; // @[Decoupled.scala 40:37]
  wire  _GEN_80; // @[LoopBlock.scala 713:33]
  wire  _GEN_81; // @[LoopBlock.scala 713:33]
  wire  _T_70; // @[Decoupled.scala 40:37]
  wire  _GEN_82; // @[LoopBlock.scala 722:57]
  wire  _GEN_83; // @[LoopBlock.scala 722:57]
  wire  _T_71; // @[Decoupled.scala 40:37]
  wire  _GEN_84; // @[LoopBlock.scala 722:57]
  wire  _GEN_85; // @[LoopBlock.scala 722:57]
  wire  _T_72; // @[Decoupled.scala 40:37]
  wire  _GEN_86; // @[LoopBlock.scala 722:57]
  wire  _GEN_87; // @[LoopBlock.scala 722:57]
  wire  _T_73; // @[Decoupled.scala 40:37]
  wire  _GEN_88; // @[LoopBlock.scala 722:57]
  wire  _GEN_89; // @[LoopBlock.scala 722:57]
  wire  _T_74; // @[Decoupled.scala 40:37]
  wire  _GEN_90; // @[LoopBlock.scala 722:57]
  wire  _GEN_91; // @[LoopBlock.scala 722:57]
  wire  _T_75; // @[Decoupled.scala 40:37]
  wire  _GEN_92; // @[LoopBlock.scala 722:57]
  wire  _GEN_93; // @[LoopBlock.scala 722:57]
  wire  _T_76; // @[Decoupled.scala 40:37]
  wire  _GEN_94; // @[LoopBlock.scala 722:57]
  wire  _GEN_95; // @[LoopBlock.scala 722:57]
  wire  _T_77; // @[Decoupled.scala 40:37]
  wire  _GEN_96; // @[LoopBlock.scala 722:57]
  wire  _GEN_97; // @[LoopBlock.scala 722:57]
  wire  _T_78; // @[Decoupled.scala 40:37]
  wire  _GEN_98; // @[LoopBlock.scala 722:57]
  wire  _GEN_99; // @[LoopBlock.scala 722:57]
  wire  _T_79; // @[Decoupled.scala 40:37]
  wire  _GEN_100; // @[LoopBlock.scala 722:57]
  wire  _GEN_101; // @[LoopBlock.scala 722:57]
  wire  _T_80; // @[Decoupled.scala 40:37]
  wire  _GEN_102; // @[LoopBlock.scala 722:57]
  wire  _GEN_103; // @[LoopBlock.scala 722:57]
  wire  _T_81; // @[Decoupled.scala 40:37]
  wire  _GEN_104; // @[LoopBlock.scala 722:57]
  wire  _GEN_105; // @[LoopBlock.scala 722:57]
  wire  _T_82; // @[Decoupled.scala 40:37]
  wire  _GEN_106; // @[LoopBlock.scala 722:57]
  wire  _GEN_107; // @[LoopBlock.scala 722:57]
  wire  _T_83; // @[Decoupled.scala 40:37]
  wire  _GEN_108; // @[LoopBlock.scala 722:57]
  wire  _GEN_109; // @[LoopBlock.scala 722:57]
  wire  _T_84; // @[Decoupled.scala 40:37]
  wire  _GEN_110; // @[LoopBlock.scala 722:57]
  wire  _GEN_111; // @[LoopBlock.scala 722:57]
  wire  _T_85; // @[Decoupled.scala 40:37]
  wire  _GEN_112; // @[LoopBlock.scala 722:57]
  wire  _GEN_113; // @[LoopBlock.scala 722:57]
  wire  _T_86; // @[Decoupled.scala 40:37]
  wire  _GEN_114; // @[LoopBlock.scala 722:57]
  wire  _GEN_115; // @[LoopBlock.scala 722:57]
  wire  _T_87; // @[Decoupled.scala 40:37]
  wire  _GEN_116; // @[LoopBlock.scala 722:57]
  wire  _GEN_117; // @[LoopBlock.scala 722:57]
  wire  _T_88; // @[Decoupled.scala 40:37]
  wire  _GEN_118; // @[LoopBlock.scala 722:57]
  wire  _GEN_119; // @[LoopBlock.scala 722:57]
  wire  _T_89; // @[Decoupled.scala 40:37]
  wire  _GEN_120; // @[LoopBlock.scala 722:57]
  wire  _GEN_121; // @[LoopBlock.scala 722:57]
  wire  _T_90; // @[Decoupled.scala 40:37]
  wire  _GEN_122; // @[LoopBlock.scala 722:57]
  wire  _GEN_123; // @[LoopBlock.scala 722:57]
  wire  _T_91; // @[Decoupled.scala 40:37]
  wire  _GEN_124; // @[LoopBlock.scala 722:57]
  wire  _GEN_125; // @[LoopBlock.scala 722:57]
  wire  _T_92; // @[Decoupled.scala 40:37]
  wire  _GEN_126; // @[LoopBlock.scala 722:57]
  wire  _GEN_127; // @[LoopBlock.scala 722:57]
  wire  _T_93; // @[Decoupled.scala 40:37]
  wire  _GEN_128; // @[LoopBlock.scala 722:57]
  wire  _GEN_129; // @[LoopBlock.scala 722:57]
  wire  _T_94; // @[Decoupled.scala 40:37]
  wire  _GEN_130; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_123;
  wire  _T_95; // @[Conditional.scala 37:30]
  wire  _T_96; // @[LoopBlock.scala 765:35]
  wire  _T_97; // @[LoopBlock.scala 765:35]
  wire  _T_98; // @[LoopBlock.scala 765:35]
  wire  _T_99; // @[LoopBlock.scala 765:35]
  wire  _T_100; // @[LoopBlock.scala 765:35]
  wire  _T_101; // @[LoopBlock.scala 765:35]
  wire  _T_102; // @[LoopBlock.scala 765:35]
  wire  _T_103; // @[LoopBlock.scala 765:35]
  wire  _T_104; // @[LoopBlock.scala 765:35]
  wire  _T_105; // @[LoopBlock.scala 765:35]
  wire  _T_106; // @[LoopBlock.scala 765:35]
  wire  _T_107; // @[LoopBlock.scala 765:35]
  wire  _T_108; // @[LoopBlock.scala 765:35]
  wire  _T_109; // @[LoopBlock.scala 765:35]
  wire  _T_110; // @[LoopBlock.scala 765:35]
  wire  _T_111; // @[LoopBlock.scala 869:28]
  wire  _GEN_132; // @[LoopBlock.scala 870:26]
  wire  _GEN_133; // @[LoopBlock.scala 870:26]
  wire  _GEN_134; // @[LoopBlock.scala 870:26]
  wire  _GEN_135; // @[LoopBlock.scala 870:26]
  wire  _GEN_136; // @[LoopBlock.scala 870:26]
  wire  _GEN_137; // @[LoopBlock.scala 870:26]
  wire  _GEN_138; // @[LoopBlock.scala 870:26]
  wire  _GEN_139; // @[LoopBlock.scala 870:26]
  wire  _GEN_140; // @[LoopBlock.scala 870:26]
  wire  _GEN_141; // @[LoopBlock.scala 870:26]
  wire  _GEN_142; // @[LoopBlock.scala 870:26]
  wire  _GEN_143; // @[LoopBlock.scala 870:26]
  wire  _GEN_144; // @[LoopBlock.scala 870:26]
  wire  _GEN_145; // @[LoopBlock.scala 870:26]
  wire  _GEN_146; // @[LoopBlock.scala 870:26]
  wire  _GEN_147; // @[LoopBlock.scala 870:26]
  wire  _GEN_148; // @[LoopBlock.scala 870:26]
  wire  _GEN_149; // @[LoopBlock.scala 870:26]
  wire  _GEN_150; // @[LoopBlock.scala 870:26]
  wire  _GEN_151; // @[LoopBlock.scala 870:26]
  wire  _GEN_152; // @[LoopBlock.scala 870:26]
  wire  _GEN_153; // @[LoopBlock.scala 870:26]
  wire  _GEN_154; // @[LoopBlock.scala 870:26]
  wire  _GEN_155; // @[LoopBlock.scala 870:26]
  wire  _GEN_156; // @[LoopBlock.scala 870:26]
  wire  _GEN_157; // @[LoopBlock.scala 870:26]
  wire  _GEN_159; // @[LoopBlock.scala 870:26]
  wire  _GEN_162; // @[LoopBlock.scala 870:26]
  wire  _GEN_164; // @[LoopBlock.scala 870:26]
  wire  _T_115; // @[Conditional.scala 37:30]
  wire  _T_116; // @[LoopBlock.scala 898:30]
  wire  _T_118; // @[LoopBlock.scala 825:65]
  wire  _T_119; // @[LoopBlock.scala 825:65]
  wire  _T_120; // @[LoopBlock.scala 825:65]
  wire  _T_121; // @[LoopBlock.scala 825:65]
  wire  _T_122; // @[LoopBlock.scala 825:65]
  wire  _T_123; // @[LoopBlock.scala 825:65]
  wire  _T_124; // @[LoopBlock.scala 825:65]
  wire  _T_125; // @[LoopBlock.scala 825:65]
  wire  _T_126; // @[LoopBlock.scala 828:26]
  wire  _T_127; // @[LoopBlock.scala 828:26]
  wire  _T_128; // @[LoopBlock.scala 828:26]
  wire  _T_129; // @[LoopBlock.scala 828:26]
  wire  _T_130; // @[LoopBlock.scala 828:26]
  wire  _T_131; // @[LoopBlock.scala 828:26]
  wire  _T_132; // @[LoopBlock.scala 828:26]
  wire  _T_133; // @[LoopBlock.scala 828:26]
  wire  _T_134; // @[LoopBlock.scala 828:26]
  wire  _T_135; // @[LoopBlock.scala 828:26]
  wire  _T_136; // @[LoopBlock.scala 828:26]
  wire  _T_137; // @[LoopBlock.scala 828:26]
  wire  _T_138; // @[LoopBlock.scala 828:26]
  wire  _T_139; // @[LoopBlock.scala 828:26]
  wire  _T_140; // @[LoopBlock.scala 828:26]
  wire  _T_141; // @[LoopBlock.scala 899:29]
  wire  _T_148; // @[LoopBlock.scala 932:19]
  wire  _T_149; // @[LoopBlock.scala 932:19]
  wire  _GEN_202; // @[LoopBlock.scala 936:64]
  wire  _GEN_205; // @[LoopBlock.scala 936:64]
  wire  _GEN_207; // @[LoopBlock.scala 936:64]
  wire  _GEN_212; // @[LoopBlock.scala 903:56]
  wire  _GEN_213; // @[LoopBlock.scala 903:56]
  wire  _GEN_215; // @[LoopBlock.scala 903:56]
  wire  _GEN_241; // @[LoopBlock.scala 903:56]
  wire  _GEN_242; // @[LoopBlock.scala 903:56]
  wire  _GEN_243; // @[LoopBlock.scala 903:56]
  wire  _GEN_244; // @[LoopBlock.scala 903:56]
  wire  _GEN_245; // @[LoopBlock.scala 903:56]
  wire  _GEN_246; // @[LoopBlock.scala 903:56]
  wire  _GEN_247; // @[LoopBlock.scala 903:56]
  wire  _GEN_248; // @[LoopBlock.scala 903:56]
  wire  _GEN_249; // @[LoopBlock.scala 903:56]
  wire  _GEN_250; // @[LoopBlock.scala 903:56]
  wire  _GEN_251; // @[LoopBlock.scala 903:56]
  wire  _GEN_252; // @[LoopBlock.scala 903:56]
  wire  _GEN_253; // @[LoopBlock.scala 903:56]
  wire  _GEN_254; // @[LoopBlock.scala 903:56]
  wire  _GEN_255; // @[LoopBlock.scala 903:56]
  wire  _GEN_256; // @[LoopBlock.scala 903:56]
  wire  _GEN_257; // @[LoopBlock.scala 903:56]
  wire  _GEN_258; // @[LoopBlock.scala 903:56]
  wire  _GEN_259; // @[LoopBlock.scala 903:56]
  wire  _GEN_260; // @[LoopBlock.scala 903:56]
  wire  _GEN_261; // @[LoopBlock.scala 903:56]
  wire  _GEN_262; // @[LoopBlock.scala 903:56]
  wire  _GEN_263; // @[LoopBlock.scala 903:56]
  wire  _GEN_264; // @[LoopBlock.scala 903:56]
  wire  _GEN_265; // @[LoopBlock.scala 903:56]
  wire  _T_157; // @[Conditional.scala 37:30]
  wire  _GEN_762; // @[LoopBlock.scala 932:19]
  wire  _GEN_763; // @[LoopBlock.scala 932:19]
  wire  _GEN_764; // @[LoopBlock.scala 932:19]
  wire  _GEN_765; // @[LoopBlock.scala 932:19]
  wire  _GEN_769; // @[LoopBlock.scala 950:19]
  wire  _GEN_770; // @[LoopBlock.scala 950:19]
  wire  _GEN_771; // @[LoopBlock.scala 950:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_28 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_28 | enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_30 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_30 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_30 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_30 | loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_32 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_32 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_32 | loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_34 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_34 | in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_36 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_36 | in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_38 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_38 | in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_40 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_40 | in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_42 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_42 | in_live_in_valid_R_4; // @[LoopBlock.scala 623:33]
  assign _T_44 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_44 | in_live_in_valid_R_5; // @[LoopBlock.scala 623:33]
  assign _T_46 = io_InLiveIn_6_ready & io_InLiveIn_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_37 = _T_46 | in_live_in_valid_R_6; // @[LoopBlock.scala 623:33]
  assign _T_48 = io_InLiveIn_7_ready & io_InLiveIn_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_41 = _T_48 | in_live_in_valid_R_7; // @[LoopBlock.scala 623:33]
  assign _T_50 = io_InLiveIn_8_ready & io_InLiveIn_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_45 = _T_50 | in_live_in_valid_R_8; // @[LoopBlock.scala 623:33]
  assign _T_52 = io_InLiveIn_9_ready & io_InLiveIn_9_valid; // @[Decoupled.scala 40:37]
  assign _GEN_49 = _T_52 | in_live_in_valid_R_9; // @[LoopBlock.scala 623:33]
  assign _T_54 = io_InLiveIn_10_ready & io_InLiveIn_10_valid; // @[Decoupled.scala 40:37]
  assign _GEN_53 = _T_54 | in_live_in_valid_R_10; // @[LoopBlock.scala 623:33]
  assign _T_56 = io_InLiveIn_11_ready & io_InLiveIn_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_57 = _T_56 | in_live_in_valid_R_11; // @[LoopBlock.scala 623:33]
  assign _T_58 = io_InLiveIn_12_ready & io_InLiveIn_12_valid; // @[Decoupled.scala 40:37]
  assign _GEN_61 = _T_58 | in_live_in_valid_R_12; // @[LoopBlock.scala 623:33]
  assign _T_60 = io_InLiveIn_13_ready & io_InLiveIn_13_valid; // @[Decoupled.scala 40:37]
  assign _GEN_65 = _T_60 | in_live_in_valid_R_13; // @[LoopBlock.scala 623:33]
  assign _T_62 = io_InLiveIn_14_ready & io_InLiveIn_14_valid; // @[Decoupled.scala 40:37]
  assign _GEN_69 = _T_62 | in_live_in_valid_R_14; // @[LoopBlock.scala 623:33]
  assign _T_64 = io_InLiveIn_15_ready & io_InLiveIn_15_valid; // @[Decoupled.scala 40:37]
  assign _GEN_73 = _T_64 | in_live_in_valid_R_15; // @[LoopBlock.scala 623:33]
  assign _T_66 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_77 = _T_66 | in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_67 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  assign _GEN_78 = _T_67 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_68 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  assign _GEN_79 = _T_68 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_69 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_80 = _T_69 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_81 = _T_69 | loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_70 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_82 = _T_70 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_83 = _T_70 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_71 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_84 = _T_71 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_85 = _T_71 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_72 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_86 = _T_72 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_87 = _T_72 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_73 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_88 = _T_73 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_89 = _T_73 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_74 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_90 = _T_74 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 722:57]
  assign _GEN_91 = _T_74 | out_live_in_fire_R_4_0; // @[LoopBlock.scala 722:57]
  assign _T_75 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_92 = _T_75 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 722:57]
  assign _GEN_93 = _T_75 | out_live_in_fire_R_5_0; // @[LoopBlock.scala 722:57]
  assign _T_76 = io_OutLiveIn_field6_0_ready & io_OutLiveIn_field6_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_94 = _T_76 ? 1'h0 : out_live_in_valid_R_6_0; // @[LoopBlock.scala 722:57]
  assign _GEN_95 = _T_76 | out_live_in_fire_R_6_0; // @[LoopBlock.scala 722:57]
  assign _T_77 = io_OutLiveIn_field7_0_ready & io_OutLiveIn_field7_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_96 = _T_77 ? 1'h0 : out_live_in_valid_R_7_0; // @[LoopBlock.scala 722:57]
  assign _GEN_97 = _T_77 | out_live_in_fire_R_7_0; // @[LoopBlock.scala 722:57]
  assign _T_78 = io_OutLiveIn_field8_0_ready & io_OutLiveIn_field8_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_98 = _T_78 ? 1'h0 : out_live_in_valid_R_8_0; // @[LoopBlock.scala 722:57]
  assign _GEN_99 = _T_78 | out_live_in_fire_R_8_0; // @[LoopBlock.scala 722:57]
  assign _T_79 = io_OutLiveIn_field9_0_ready & io_OutLiveIn_field9_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_100 = _T_79 ? 1'h0 : out_live_in_valid_R_9_0; // @[LoopBlock.scala 722:57]
  assign _GEN_101 = _T_79 | out_live_in_fire_R_9_0; // @[LoopBlock.scala 722:57]
  assign _T_80 = io_OutLiveIn_field10_0_ready & io_OutLiveIn_field10_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_102 = _T_80 ? 1'h0 : out_live_in_valid_R_10_0; // @[LoopBlock.scala 722:57]
  assign _GEN_103 = _T_80 | out_live_in_fire_R_10_0; // @[LoopBlock.scala 722:57]
  assign _T_81 = io_OutLiveIn_field10_1_ready & io_OutLiveIn_field10_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_104 = _T_81 ? 1'h0 : out_live_in_valid_R_10_1; // @[LoopBlock.scala 722:57]
  assign _GEN_105 = _T_81 | out_live_in_fire_R_10_1; // @[LoopBlock.scala 722:57]
  assign _T_82 = io_OutLiveIn_field10_2_ready & io_OutLiveIn_field10_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_106 = _T_82 ? 1'h0 : out_live_in_valid_R_10_2; // @[LoopBlock.scala 722:57]
  assign _GEN_107 = _T_82 | out_live_in_fire_R_10_2; // @[LoopBlock.scala 722:57]
  assign _T_83 = io_OutLiveIn_field10_3_ready & io_OutLiveIn_field10_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_108 = _T_83 ? 1'h0 : out_live_in_valid_R_10_3; // @[LoopBlock.scala 722:57]
  assign _GEN_109 = _T_83 | out_live_in_fire_R_10_3; // @[LoopBlock.scala 722:57]
  assign _T_84 = io_OutLiveIn_field10_4_ready & io_OutLiveIn_field10_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_110 = _T_84 ? 1'h0 : out_live_in_valid_R_10_4; // @[LoopBlock.scala 722:57]
  assign _GEN_111 = _T_84 | out_live_in_fire_R_10_4; // @[LoopBlock.scala 722:57]
  assign _T_85 = io_OutLiveIn_field10_5_ready & io_OutLiveIn_field10_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_112 = _T_85 ? 1'h0 : out_live_in_valid_R_10_5; // @[LoopBlock.scala 722:57]
  assign _GEN_113 = _T_85 | out_live_in_fire_R_10_5; // @[LoopBlock.scala 722:57]
  assign _T_86 = io_OutLiveIn_field10_6_ready & io_OutLiveIn_field10_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_114 = _T_86 ? 1'h0 : out_live_in_valid_R_10_6; // @[LoopBlock.scala 722:57]
  assign _GEN_115 = _T_86 | out_live_in_fire_R_10_6; // @[LoopBlock.scala 722:57]
  assign _T_87 = io_OutLiveIn_field10_7_ready & io_OutLiveIn_field10_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_116 = _T_87 ? 1'h0 : out_live_in_valid_R_10_7; // @[LoopBlock.scala 722:57]
  assign _GEN_117 = _T_87 | out_live_in_fire_R_10_7; // @[LoopBlock.scala 722:57]
  assign _T_88 = io_OutLiveIn_field10_8_ready & io_OutLiveIn_field10_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_118 = _T_88 ? 1'h0 : out_live_in_valid_R_10_8; // @[LoopBlock.scala 722:57]
  assign _GEN_119 = _T_88 | out_live_in_fire_R_10_8; // @[LoopBlock.scala 722:57]
  assign _T_89 = io_OutLiveIn_field11_0_ready & io_OutLiveIn_field11_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_120 = _T_89 ? 1'h0 : out_live_in_valid_R_11_0; // @[LoopBlock.scala 722:57]
  assign _GEN_121 = _T_89 | out_live_in_fire_R_11_0; // @[LoopBlock.scala 722:57]
  assign _T_90 = io_OutLiveIn_field12_0_ready & io_OutLiveIn_field12_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_122 = _T_90 ? 1'h0 : out_live_in_valid_R_12_0; // @[LoopBlock.scala 722:57]
  assign _GEN_123 = _T_90 | out_live_in_fire_R_12_0; // @[LoopBlock.scala 722:57]
  assign _T_91 = io_OutLiveIn_field13_0_ready & io_OutLiveIn_field13_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_124 = _T_91 ? 1'h0 : out_live_in_valid_R_13_0; // @[LoopBlock.scala 722:57]
  assign _GEN_125 = _T_91 | out_live_in_fire_R_13_0; // @[LoopBlock.scala 722:57]
  assign _T_92 = io_OutLiveIn_field14_0_ready & io_OutLiveIn_field14_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_126 = _T_92 ? 1'h0 : out_live_in_valid_R_14_0; // @[LoopBlock.scala 722:57]
  assign _GEN_127 = _T_92 | out_live_in_fire_R_14_0; // @[LoopBlock.scala 722:57]
  assign _T_93 = io_OutLiveIn_field15_0_ready & io_OutLiveIn_field15_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_128 = _T_93 ? 1'h0 : out_live_in_valid_R_15_0; // @[LoopBlock.scala 722:57]
  assign _GEN_129 = _T_93 | out_live_in_fire_R_15_0; // @[LoopBlock.scala 722:57]
  assign _T_94 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_130 = _T_94 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_95 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_96 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_97 = _T_96 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_98 = _T_97 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_99 = _T_98 & in_live_in_valid_R_4; // @[LoopBlock.scala 765:35]
  assign _T_100 = _T_99 & in_live_in_valid_R_5; // @[LoopBlock.scala 765:35]
  assign _T_101 = _T_100 & in_live_in_valid_R_6; // @[LoopBlock.scala 765:35]
  assign _T_102 = _T_101 & in_live_in_valid_R_7; // @[LoopBlock.scala 765:35]
  assign _T_103 = _T_102 & in_live_in_valid_R_8; // @[LoopBlock.scala 765:35]
  assign _T_104 = _T_103 & in_live_in_valid_R_9; // @[LoopBlock.scala 765:35]
  assign _T_105 = _T_104 & in_live_in_valid_R_10; // @[LoopBlock.scala 765:35]
  assign _T_106 = _T_105 & in_live_in_valid_R_11; // @[LoopBlock.scala 765:35]
  assign _T_107 = _T_106 & in_live_in_valid_R_12; // @[LoopBlock.scala 765:35]
  assign _T_108 = _T_107 & in_live_in_valid_R_13; // @[LoopBlock.scala 765:35]
  assign _T_109 = _T_108 & in_live_in_valid_R_14; // @[LoopBlock.scala 765:35]
  assign _T_110 = _T_109 & in_live_in_valid_R_15; // @[LoopBlock.scala 765:35]
  assign _T_111 = _T_110 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_132 = enable_R_control | _GEN_82; // @[LoopBlock.scala 870:26]
  assign _GEN_133 = enable_R_control | _GEN_84; // @[LoopBlock.scala 870:26]
  assign _GEN_134 = enable_R_control | _GEN_86; // @[LoopBlock.scala 870:26]
  assign _GEN_135 = enable_R_control | _GEN_88; // @[LoopBlock.scala 870:26]
  assign _GEN_136 = enable_R_control | _GEN_90; // @[LoopBlock.scala 870:26]
  assign _GEN_137 = enable_R_control | _GEN_92; // @[LoopBlock.scala 870:26]
  assign _GEN_138 = enable_R_control | _GEN_94; // @[LoopBlock.scala 870:26]
  assign _GEN_139 = enable_R_control | _GEN_96; // @[LoopBlock.scala 870:26]
  assign _GEN_140 = enable_R_control | _GEN_98; // @[LoopBlock.scala 870:26]
  assign _GEN_141 = enable_R_control | _GEN_100; // @[LoopBlock.scala 870:26]
  assign _GEN_142 = enable_R_control | _GEN_102; // @[LoopBlock.scala 870:26]
  assign _GEN_143 = enable_R_control | _GEN_104; // @[LoopBlock.scala 870:26]
  assign _GEN_144 = enable_R_control | _GEN_106; // @[LoopBlock.scala 870:26]
  assign _GEN_145 = enable_R_control | _GEN_108; // @[LoopBlock.scala 870:26]
  assign _GEN_146 = enable_R_control | _GEN_110; // @[LoopBlock.scala 870:26]
  assign _GEN_147 = enable_R_control | _GEN_112; // @[LoopBlock.scala 870:26]
  assign _GEN_148 = enable_R_control | _GEN_114; // @[LoopBlock.scala 870:26]
  assign _GEN_149 = enable_R_control | _GEN_116; // @[LoopBlock.scala 870:26]
  assign _GEN_150 = enable_R_control | _GEN_118; // @[LoopBlock.scala 870:26]
  assign _GEN_151 = enable_R_control | _GEN_120; // @[LoopBlock.scala 870:26]
  assign _GEN_152 = enable_R_control | _GEN_122; // @[LoopBlock.scala 870:26]
  assign _GEN_153 = enable_R_control | _GEN_124; // @[LoopBlock.scala 870:26]
  assign _GEN_154 = enable_R_control | _GEN_126; // @[LoopBlock.scala 870:26]
  assign _GEN_155 = enable_R_control | _GEN_128; // @[LoopBlock.scala 870:26]
  assign _GEN_156 = enable_R_control | _GEN_130; // @[LoopBlock.scala 870:26]
  assign _GEN_157 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_159 = enable_R_control | _GEN_78; // @[LoopBlock.scala 870:26]
  assign _GEN_162 = enable_R_control | _GEN_79; // @[LoopBlock.scala 870:26]
  assign _GEN_164 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 870:26]
  assign _T_115 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_116 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_118 = out_live_in_fire_R_10_0 & out_live_in_fire_R_10_1; // @[LoopBlock.scala 825:65]
  assign _T_119 = _T_118 & out_live_in_fire_R_10_2; // @[LoopBlock.scala 825:65]
  assign _T_120 = _T_119 & out_live_in_fire_R_10_3; // @[LoopBlock.scala 825:65]
  assign _T_121 = _T_120 & out_live_in_fire_R_10_4; // @[LoopBlock.scala 825:65]
  assign _T_122 = _T_121 & out_live_in_fire_R_10_5; // @[LoopBlock.scala 825:65]
  assign _T_123 = _T_122 & out_live_in_fire_R_10_6; // @[LoopBlock.scala 825:65]
  assign _T_124 = _T_123 & out_live_in_fire_R_10_7; // @[LoopBlock.scala 825:65]
  assign _T_125 = _T_124 & out_live_in_fire_R_10_8; // @[LoopBlock.scala 825:65]
  assign _T_126 = out_live_in_fire_R_0_0 & out_live_in_fire_R_1_0; // @[LoopBlock.scala 828:26]
  assign _T_127 = _T_126 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_128 = _T_127 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_129 = _T_128 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 828:26]
  assign _T_130 = _T_129 & out_live_in_fire_R_5_0; // @[LoopBlock.scala 828:26]
  assign _T_131 = _T_130 & out_live_in_fire_R_6_0; // @[LoopBlock.scala 828:26]
  assign _T_132 = _T_131 & out_live_in_fire_R_7_0; // @[LoopBlock.scala 828:26]
  assign _T_133 = _T_132 & out_live_in_fire_R_8_0; // @[LoopBlock.scala 828:26]
  assign _T_134 = _T_133 & out_live_in_fire_R_9_0; // @[LoopBlock.scala 828:26]
  assign _T_135 = _T_134 & _T_125; // @[LoopBlock.scala 828:26]
  assign _T_136 = _T_135 & out_live_in_fire_R_11_0; // @[LoopBlock.scala 828:26]
  assign _T_137 = _T_136 & out_live_in_fire_R_12_0; // @[LoopBlock.scala 828:26]
  assign _T_138 = _T_137 & out_live_in_fire_R_13_0; // @[LoopBlock.scala 828:26]
  assign _T_139 = _T_138 & out_live_in_fire_R_14_0; // @[LoopBlock.scala 828:26]
  assign _T_140 = _T_139 & out_live_in_fire_R_15_0; // @[LoopBlock.scala 828:26]
  assign _T_141 = _T_116 & _T_140; // @[LoopBlock.scala 899:29]
  assign _T_148 = $unsigned(reset); // @[LoopBlock.scala 932:19]
  assign _T_149 = _T_148 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_202 = loop_finish_R_0_control | _GEN_80; // @[LoopBlock.scala 936:64]
  assign _GEN_205 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_207 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_212 = loop_back_R_0_control | _GEN_78; // @[LoopBlock.scala 903:56]
  assign _GEN_213 = loop_back_R_0_control | _GEN_205; // @[LoopBlock.scala 903:56]
  assign _GEN_215 = loop_back_R_0_control | _GEN_79; // @[LoopBlock.scala 903:56]
  assign _GEN_241 = loop_back_R_0_control | _GEN_82; // @[LoopBlock.scala 903:56]
  assign _GEN_242 = loop_back_R_0_control | _GEN_84; // @[LoopBlock.scala 903:56]
  assign _GEN_243 = loop_back_R_0_control | _GEN_86; // @[LoopBlock.scala 903:56]
  assign _GEN_244 = loop_back_R_0_control | _GEN_88; // @[LoopBlock.scala 903:56]
  assign _GEN_245 = loop_back_R_0_control | _GEN_90; // @[LoopBlock.scala 903:56]
  assign _GEN_246 = loop_back_R_0_control | _GEN_92; // @[LoopBlock.scala 903:56]
  assign _GEN_247 = loop_back_R_0_control | _GEN_94; // @[LoopBlock.scala 903:56]
  assign _GEN_248 = loop_back_R_0_control | _GEN_96; // @[LoopBlock.scala 903:56]
  assign _GEN_249 = loop_back_R_0_control | _GEN_98; // @[LoopBlock.scala 903:56]
  assign _GEN_250 = loop_back_R_0_control | _GEN_100; // @[LoopBlock.scala 903:56]
  assign _GEN_251 = loop_back_R_0_control | _GEN_102; // @[LoopBlock.scala 903:56]
  assign _GEN_252 = loop_back_R_0_control | _GEN_104; // @[LoopBlock.scala 903:56]
  assign _GEN_253 = loop_back_R_0_control | _GEN_106; // @[LoopBlock.scala 903:56]
  assign _GEN_254 = loop_back_R_0_control | _GEN_108; // @[LoopBlock.scala 903:56]
  assign _GEN_255 = loop_back_R_0_control | _GEN_110; // @[LoopBlock.scala 903:56]
  assign _GEN_256 = loop_back_R_0_control | _GEN_112; // @[LoopBlock.scala 903:56]
  assign _GEN_257 = loop_back_R_0_control | _GEN_114; // @[LoopBlock.scala 903:56]
  assign _GEN_258 = loop_back_R_0_control | _GEN_116; // @[LoopBlock.scala 903:56]
  assign _GEN_259 = loop_back_R_0_control | _GEN_118; // @[LoopBlock.scala 903:56]
  assign _GEN_260 = loop_back_R_0_control | _GEN_120; // @[LoopBlock.scala 903:56]
  assign _GEN_261 = loop_back_R_0_control | _GEN_122; // @[LoopBlock.scala 903:56]
  assign _GEN_262 = loop_back_R_0_control | _GEN_124; // @[LoopBlock.scala 903:56]
  assign _GEN_263 = loop_back_R_0_control | _GEN_126; // @[LoopBlock.scala 903:56]
  assign _GEN_264 = loop_back_R_0_control | _GEN_128; // @[LoopBlock.scala 903:56]
  assign _GEN_265 = loop_back_R_0_control | _GEN_130; // @[LoopBlock.scala 903:56]
  assign _T_157 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_4_ready = ~ in_live_in_valid_R_4; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_5_ready = ~ in_live_in_valid_R_5; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_6_ready = ~ in_live_in_valid_R_6; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_7_ready = ~ in_live_in_valid_R_7; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_8_ready = ~ in_live_in_valid_R_8; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_9_ready = ~ in_live_in_valid_R_9; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_10_ready = ~ in_live_in_valid_R_10; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_11_ready = ~ in_live_in_valid_R_11; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_12_ready = ~ in_live_in_valid_R_12; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_13_ready = ~ in_live_in_valid_R_13; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_14_ready = ~ in_live_in_valid_R_14; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_15_ready = ~ in_live_in_valid_R_15; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field15_0_valid = out_live_in_valid_R_15_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field15_0_bits_predicate = in_live_in_R_15_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field15_0_bits_taskID = in_live_in_R_15_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field15_0_bits_data = in_live_in_R_15_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field14_0_valid = out_live_in_valid_R_14_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field14_0_bits_predicate = in_live_in_R_14_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field14_0_bits_taskID = in_live_in_R_14_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field14_0_bits_data = in_live_in_R_14_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field13_0_valid = out_live_in_valid_R_13_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field13_0_bits_predicate = in_live_in_R_13_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field13_0_bits_taskID = in_live_in_R_13_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field13_0_bits_data = in_live_in_R_13_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field12_0_valid = out_live_in_valid_R_12_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field12_0_bits_predicate = in_live_in_R_12_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field12_0_bits_taskID = in_live_in_R_12_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field12_0_bits_data = in_live_in_R_12_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field11_0_valid = out_live_in_valid_R_11_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field11_0_bits_taskID = in_live_in_R_11_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field11_0_bits_data = in_live_in_R_11_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_0_valid = out_live_in_valid_R_10_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_0_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_0_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_1_valid = out_live_in_valid_R_10_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_1_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_1_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_2_valid = out_live_in_valid_R_10_2; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_2_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_2_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_3_valid = out_live_in_valid_R_10_3; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_3_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_3_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_4_valid = out_live_in_valid_R_10_4; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_4_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_4_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_5_valid = out_live_in_valid_R_10_5; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_5_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_5_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_6_valid = out_live_in_valid_R_10_6; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_6_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_6_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_7_valid = out_live_in_valid_R_10_7; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_7_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_7_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_8_valid = out_live_in_valid_R_10_8; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_8_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_8_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field9_0_valid = out_live_in_valid_R_9_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field9_0_bits_predicate = in_live_in_R_9_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field9_0_bits_taskID = in_live_in_R_9_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field9_0_bits_data = in_live_in_R_9_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_valid = out_live_in_valid_R_8_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field8_0_bits_predicate = in_live_in_R_8_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_bits_taskID = in_live_in_R_8_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_bits_data = in_live_in_R_8_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_valid = out_live_in_valid_R_7_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field7_0_bits_predicate = in_live_in_R_7_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_bits_taskID = in_live_in_R_7_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_bits_data = in_live_in_R_7_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_valid = out_live_in_valid_R_6_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field6_0_bits_predicate = in_live_in_R_6_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_bits_taskID = in_live_in_R_6_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_bits_data = in_live_in_R_6_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_0_bits_predicate = in_live_in_R_4_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_bits_taskID = in_live_in_R_4_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
  assign _GEN_762 = _T_95 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_763 = _GEN_762 & _T_115; // @[LoopBlock.scala 932:19]
  assign _GEN_764 = _GEN_763 & _T_141; // @[LoopBlock.scala 932:19]
  assign _GEN_765 = _GEN_764 & loop_back_R_0_control; // @[LoopBlock.scala 932:19]
  assign _GEN_769 = loop_back_R_0_control == 1'h0; // @[LoopBlock.scala 950:19]
  assign _GEN_770 = _GEN_764 & _GEN_769; // @[LoopBlock.scala 950:19]
  assign _GEN_771 = _GEN_770 & loop_finish_R_0_control; // @[LoopBlock.scala 950:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_4_predicate = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_4_taskID = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_R_4_data = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_R_5_data = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_R_6_predicate = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_R_6_taskID = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_live_in_R_6_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_live_in_R_7_predicate = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_live_in_R_7_taskID = _RAND_21[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_live_in_R_7_data = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_live_in_R_8_predicate = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_live_in_R_8_taskID = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_live_in_R_8_data = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  in_live_in_R_9_predicate = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  in_live_in_R_9_taskID = _RAND_27[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  in_live_in_R_9_data = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  in_live_in_R_10_taskID = _RAND_29[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  in_live_in_R_10_data = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  in_live_in_R_11_taskID = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  in_live_in_R_11_data = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  in_live_in_R_12_predicate = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  in_live_in_R_12_taskID = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  in_live_in_R_12_data = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  in_live_in_R_13_predicate = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  in_live_in_R_13_taskID = _RAND_37[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  in_live_in_R_13_data = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  in_live_in_R_14_predicate = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  in_live_in_R_14_taskID = _RAND_40[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  in_live_in_R_14_data = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  in_live_in_R_15_predicate = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  in_live_in_R_15_taskID = _RAND_43[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  in_live_in_R_15_data = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  in_live_in_valid_R_6 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  in_live_in_valid_R_7 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  in_live_in_valid_R_8 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  in_live_in_valid_R_9 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  in_live_in_valid_R_10 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  in_live_in_valid_R_11 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  in_live_in_valid_R_12 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  in_live_in_valid_R_13 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  in_live_in_valid_R_14 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  in_live_in_valid_R_15 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_61[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  out_live_in_valid_R_6_0 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  out_live_in_valid_R_7_0 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  out_live_in_valid_R_8_0 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  out_live_in_valid_R_9_0 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  out_live_in_valid_R_10_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  out_live_in_valid_R_10_1 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  out_live_in_valid_R_10_2 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  out_live_in_valid_R_10_3 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  out_live_in_valid_R_10_4 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  out_live_in_valid_R_10_5 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  out_live_in_valid_R_10_6 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  out_live_in_valid_R_10_7 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  out_live_in_valid_R_10_8 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  out_live_in_valid_R_11_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  out_live_in_valid_R_12_0 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  out_live_in_valid_R_13_0 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  out_live_in_valid_R_14_0 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  out_live_in_valid_R_15_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  out_live_in_fire_R_6_0 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  out_live_in_fire_R_7_0 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  out_live_in_fire_R_8_0 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  out_live_in_fire_R_9_0 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  out_live_in_fire_R_10_0 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  out_live_in_fire_R_10_1 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  out_live_in_fire_R_10_2 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  out_live_in_fire_R_10_3 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  out_live_in_fire_R_10_4 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  out_live_in_fire_R_10_5 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  out_live_in_fire_R_10_6 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  out_live_in_fire_R_10_7 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  out_live_in_fire_R_10_8 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  out_live_in_fire_R_11_0 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  out_live_in_fire_R_12_0 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  out_live_in_fire_R_13_0 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  out_live_in_fire_R_14_0 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  out_live_in_fire_R_15_0 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_113[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_116[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_119[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  state = _RAND_123[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_28) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_28) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_28) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_28) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_28) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_115) begin
          if (_T_28) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_28) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_28) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_95) begin
        enable_valid_R <= _GEN_3;
      end else begin
        if (_T_115) begin
          enable_valid_R <= _GEN_3;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_3;
            end
          end else begin
            enable_valid_R <= _GEN_3;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_30) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_30) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_30) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_30) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_30) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_30) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_30) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_30) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        loop_back_valid_R_0 <= _GEN_6;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_32) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_32) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_32) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_32) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_7;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        loop_finish_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_34) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_34) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_34) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_34) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_36) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_36) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_36) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_36) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_38) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_38) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_38) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_38) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_40) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_40) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_40) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_40) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_predicate <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_42) begin
          in_live_in_R_4_predicate <= io_InLiveIn_4_bits_predicate;
        end
      end else begin
        if (_T_115) begin
          if (_T_42) begin
            in_live_in_R_4_predicate <= io_InLiveIn_4_bits_predicate;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_predicate <= 1'h0;
            end else begin
              if (_T_42) begin
                in_live_in_R_4_predicate <= io_InLiveIn_4_bits_predicate;
              end
            end
          end else begin
            if (_T_42) begin
              in_live_in_R_4_predicate <= io_InLiveIn_4_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_42) begin
          in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_42) begin
            in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_taskID <= 5'h0;
            end else begin
              if (_T_42) begin
                in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
              end
            end
          end else begin
            if (_T_42) begin
              in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_42) begin
          in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_42) begin
            in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_data <= 32'h0;
            end else begin
              if (_T_42) begin
                in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
              end
            end
          end else begin
            if (_T_42) begin
              in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_44) begin
          in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_44) begin
            in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_data <= 32'h0;
            end else begin
              if (_T_44) begin
                in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
              end
            end
          end else begin
            if (_T_44) begin
              in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_predicate <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_46) begin
          in_live_in_R_6_predicate <= io_InLiveIn_6_bits_predicate;
        end
      end else begin
        if (_T_115) begin
          if (_T_46) begin
            in_live_in_R_6_predicate <= io_InLiveIn_6_bits_predicate;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_predicate <= 1'h0;
            end else begin
              if (_T_46) begin
                in_live_in_R_6_predicate <= io_InLiveIn_6_bits_predicate;
              end
            end
          end else begin
            if (_T_46) begin
              in_live_in_R_6_predicate <= io_InLiveIn_6_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_46) begin
          in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_46) begin
            in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_taskID <= 5'h0;
            end else begin
              if (_T_46) begin
                in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
              end
            end
          end else begin
            if (_T_46) begin
              in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_46) begin
          in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_46) begin
            in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_data <= 32'h0;
            end else begin
              if (_T_46) begin
                in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
              end
            end
          end else begin
            if (_T_46) begin
              in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_predicate <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_48) begin
          in_live_in_R_7_predicate <= io_InLiveIn_7_bits_predicate;
        end
      end else begin
        if (_T_115) begin
          if (_T_48) begin
            in_live_in_R_7_predicate <= io_InLiveIn_7_bits_predicate;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_predicate <= 1'h0;
            end else begin
              if (_T_48) begin
                in_live_in_R_7_predicate <= io_InLiveIn_7_bits_predicate;
              end
            end
          end else begin
            if (_T_48) begin
              in_live_in_R_7_predicate <= io_InLiveIn_7_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_48) begin
          in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_48) begin
            in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_taskID <= 5'h0;
            end else begin
              if (_T_48) begin
                in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
              end
            end
          end else begin
            if (_T_48) begin
              in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_48) begin
          in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_48) begin
            in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_data <= 32'h0;
            end else begin
              if (_T_48) begin
                in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
              end
            end
          end else begin
            if (_T_48) begin
              in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_predicate <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_50) begin
          in_live_in_R_8_predicate <= io_InLiveIn_8_bits_predicate;
        end
      end else begin
        if (_T_115) begin
          if (_T_50) begin
            in_live_in_R_8_predicate <= io_InLiveIn_8_bits_predicate;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_predicate <= 1'h0;
            end else begin
              if (_T_50) begin
                in_live_in_R_8_predicate <= io_InLiveIn_8_bits_predicate;
              end
            end
          end else begin
            if (_T_50) begin
              in_live_in_R_8_predicate <= io_InLiveIn_8_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_50) begin
          in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_50) begin
            in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_taskID <= 5'h0;
            end else begin
              if (_T_50) begin
                in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
              end
            end
          end else begin
            if (_T_50) begin
              in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_50) begin
          in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_50) begin
            in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_data <= 32'h0;
            end else begin
              if (_T_50) begin
                in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
              end
            end
          end else begin
            if (_T_50) begin
              in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_9_predicate <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_52) begin
          in_live_in_R_9_predicate <= io_InLiveIn_9_bits_predicate;
        end
      end else begin
        if (_T_115) begin
          if (_T_52) begin
            in_live_in_R_9_predicate <= io_InLiveIn_9_bits_predicate;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_9_predicate <= 1'h0;
            end else begin
              if (_T_52) begin
                in_live_in_R_9_predicate <= io_InLiveIn_9_bits_predicate;
              end
            end
          end else begin
            if (_T_52) begin
              in_live_in_R_9_predicate <= io_InLiveIn_9_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_9_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_52) begin
          in_live_in_R_9_taskID <= io_InLiveIn_9_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_52) begin
            in_live_in_R_9_taskID <= io_InLiveIn_9_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_9_taskID <= 5'h0;
            end else begin
              if (_T_52) begin
                in_live_in_R_9_taskID <= io_InLiveIn_9_bits_taskID;
              end
            end
          end else begin
            if (_T_52) begin
              in_live_in_R_9_taskID <= io_InLiveIn_9_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_9_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_52) begin
          in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_52) begin
            in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_9_data <= 32'h0;
            end else begin
              if (_T_52) begin
                in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
              end
            end
          end else begin
            if (_T_52) begin
              in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_10_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_54) begin
          in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_54) begin
            in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_10_taskID <= 5'h0;
            end else begin
              if (_T_54) begin
                in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
              end
            end
          end else begin
            if (_T_54) begin
              in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_10_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_54) begin
          in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_54) begin
            in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_10_data <= 32'h0;
            end else begin
              if (_T_54) begin
                in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
              end
            end
          end else begin
            if (_T_54) begin
              in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_11_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_56) begin
          in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_56) begin
            in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_11_taskID <= 5'h0;
            end else begin
              if (_T_56) begin
                in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
              end
            end
          end else begin
            if (_T_56) begin
              in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_11_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_56) begin
          in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_56) begin
            in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_11_data <= 32'h0;
            end else begin
              if (_T_56) begin
                in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
              end
            end
          end else begin
            if (_T_56) begin
              in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_12_predicate <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_58) begin
          in_live_in_R_12_predicate <= io_InLiveIn_12_bits_predicate;
        end
      end else begin
        if (_T_115) begin
          if (_T_58) begin
            in_live_in_R_12_predicate <= io_InLiveIn_12_bits_predicate;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_12_predicate <= 1'h0;
            end else begin
              if (_T_58) begin
                in_live_in_R_12_predicate <= io_InLiveIn_12_bits_predicate;
              end
            end
          end else begin
            if (_T_58) begin
              in_live_in_R_12_predicate <= io_InLiveIn_12_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_12_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_58) begin
          in_live_in_R_12_taskID <= io_InLiveIn_12_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_58) begin
            in_live_in_R_12_taskID <= io_InLiveIn_12_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_12_taskID <= 5'h0;
            end else begin
              if (_T_58) begin
                in_live_in_R_12_taskID <= io_InLiveIn_12_bits_taskID;
              end
            end
          end else begin
            if (_T_58) begin
              in_live_in_R_12_taskID <= io_InLiveIn_12_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_12_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_58) begin
          in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_58) begin
            in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_12_data <= 32'h0;
            end else begin
              if (_T_58) begin
                in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
              end
            end
          end else begin
            if (_T_58) begin
              in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_13_predicate <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_60) begin
          in_live_in_R_13_predicate <= io_InLiveIn_13_bits_predicate;
        end
      end else begin
        if (_T_115) begin
          if (_T_60) begin
            in_live_in_R_13_predicate <= io_InLiveIn_13_bits_predicate;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_13_predicate <= 1'h0;
            end else begin
              if (_T_60) begin
                in_live_in_R_13_predicate <= io_InLiveIn_13_bits_predicate;
              end
            end
          end else begin
            if (_T_60) begin
              in_live_in_R_13_predicate <= io_InLiveIn_13_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_13_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_60) begin
          in_live_in_R_13_taskID <= io_InLiveIn_13_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_60) begin
            in_live_in_R_13_taskID <= io_InLiveIn_13_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_13_taskID <= 5'h0;
            end else begin
              if (_T_60) begin
                in_live_in_R_13_taskID <= io_InLiveIn_13_bits_taskID;
              end
            end
          end else begin
            if (_T_60) begin
              in_live_in_R_13_taskID <= io_InLiveIn_13_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_13_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_60) begin
          in_live_in_R_13_data <= io_InLiveIn_13_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_60) begin
            in_live_in_R_13_data <= io_InLiveIn_13_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_13_data <= 32'h0;
            end else begin
              if (_T_60) begin
                in_live_in_R_13_data <= io_InLiveIn_13_bits_data;
              end
            end
          end else begin
            if (_T_60) begin
              in_live_in_R_13_data <= io_InLiveIn_13_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_14_predicate <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_62) begin
          in_live_in_R_14_predicate <= io_InLiveIn_14_bits_predicate;
        end
      end else begin
        if (_T_115) begin
          if (_T_62) begin
            in_live_in_R_14_predicate <= io_InLiveIn_14_bits_predicate;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_14_predicate <= 1'h0;
            end else begin
              if (_T_62) begin
                in_live_in_R_14_predicate <= io_InLiveIn_14_bits_predicate;
              end
            end
          end else begin
            if (_T_62) begin
              in_live_in_R_14_predicate <= io_InLiveIn_14_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_14_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_62) begin
          in_live_in_R_14_taskID <= io_InLiveIn_14_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_62) begin
            in_live_in_R_14_taskID <= io_InLiveIn_14_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_14_taskID <= 5'h0;
            end else begin
              if (_T_62) begin
                in_live_in_R_14_taskID <= io_InLiveIn_14_bits_taskID;
              end
            end
          end else begin
            if (_T_62) begin
              in_live_in_R_14_taskID <= io_InLiveIn_14_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_14_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_62) begin
          in_live_in_R_14_data <= io_InLiveIn_14_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_62) begin
            in_live_in_R_14_data <= io_InLiveIn_14_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_14_data <= 32'h0;
            end else begin
              if (_T_62) begin
                in_live_in_R_14_data <= io_InLiveIn_14_bits_data;
              end
            end
          end else begin
            if (_T_62) begin
              in_live_in_R_14_data <= io_InLiveIn_14_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_15_predicate <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_64) begin
          in_live_in_R_15_predicate <= io_InLiveIn_15_bits_predicate;
        end
      end else begin
        if (_T_115) begin
          if (_T_64) begin
            in_live_in_R_15_predicate <= io_InLiveIn_15_bits_predicate;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_15_predicate <= 1'h0;
            end else begin
              if (_T_64) begin
                in_live_in_R_15_predicate <= io_InLiveIn_15_bits_predicate;
              end
            end
          end else begin
            if (_T_64) begin
              in_live_in_R_15_predicate <= io_InLiveIn_15_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_15_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_64) begin
          in_live_in_R_15_taskID <= io_InLiveIn_15_bits_taskID;
        end
      end else begin
        if (_T_115) begin
          if (_T_64) begin
            in_live_in_R_15_taskID <= io_InLiveIn_15_bits_taskID;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_15_taskID <= 5'h0;
            end else begin
              if (_T_64) begin
                in_live_in_R_15_taskID <= io_InLiveIn_15_bits_taskID;
              end
            end
          end else begin
            if (_T_64) begin
              in_live_in_R_15_taskID <= io_InLiveIn_15_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_15_data <= 32'h0;
    end else begin
      if (_T_95) begin
        if (_T_64) begin
          in_live_in_R_15_data <= io_InLiveIn_15_bits_data;
        end
      end else begin
        if (_T_115) begin
          if (_T_64) begin
            in_live_in_R_15_data <= io_InLiveIn_15_bits_data;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_15_data <= 32'h0;
            end else begin
              if (_T_64) begin
                in_live_in_R_15_data <= io_InLiveIn_15_bits_data;
              end
            end
          end else begin
            if (_T_64) begin
              in_live_in_R_15_data <= io_InLiveIn_15_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_0 <= _GEN_13;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_0 <= _GEN_13;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              in_live_in_valid_R_0 <= _GEN_13;
            end
          end else begin
            in_live_in_valid_R_0 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_1 <= _GEN_17;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_1 <= _GEN_17;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              in_live_in_valid_R_1 <= _GEN_17;
            end
          end else begin
            in_live_in_valid_R_1 <= _GEN_17;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_2 <= _GEN_21;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              in_live_in_valid_R_2 <= _GEN_21;
            end
          end else begin
            in_live_in_valid_R_2 <= _GEN_21;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_3 <= _GEN_25;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_3 <= _GEN_25;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              in_live_in_valid_R_3 <= _GEN_25;
            end
          end else begin
            in_live_in_valid_R_3 <= _GEN_25;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_4 <= _GEN_29;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_4 <= _GEN_29;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_4 <= 1'h0;
            end else begin
              in_live_in_valid_R_4 <= _GEN_29;
            end
          end else begin
            in_live_in_valid_R_4 <= _GEN_29;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_5 <= _GEN_33;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_5 <= _GEN_33;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_5 <= 1'h0;
            end else begin
              in_live_in_valid_R_5 <= _GEN_33;
            end
          end else begin
            in_live_in_valid_R_5 <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_6 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_6 <= _GEN_37;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_6 <= _GEN_37;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_6 <= 1'h0;
            end else begin
              in_live_in_valid_R_6 <= _GEN_37;
            end
          end else begin
            in_live_in_valid_R_6 <= _GEN_37;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_7 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_7 <= _GEN_41;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_7 <= _GEN_41;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_7 <= 1'h0;
            end else begin
              in_live_in_valid_R_7 <= _GEN_41;
            end
          end else begin
            in_live_in_valid_R_7 <= _GEN_41;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_8 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_8 <= _GEN_45;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_8 <= _GEN_45;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_8 <= 1'h0;
            end else begin
              in_live_in_valid_R_8 <= _GEN_45;
            end
          end else begin
            in_live_in_valid_R_8 <= _GEN_45;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_9 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_9 <= _GEN_49;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_9 <= _GEN_49;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_9 <= 1'h0;
            end else begin
              in_live_in_valid_R_9 <= _GEN_49;
            end
          end else begin
            in_live_in_valid_R_9 <= _GEN_49;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_10 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_10 <= _GEN_53;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_10 <= _GEN_53;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_10 <= 1'h0;
            end else begin
              in_live_in_valid_R_10 <= _GEN_53;
            end
          end else begin
            in_live_in_valid_R_10 <= _GEN_53;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_11 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_11 <= _GEN_57;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_11 <= _GEN_57;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_11 <= 1'h0;
            end else begin
              in_live_in_valid_R_11 <= _GEN_57;
            end
          end else begin
            in_live_in_valid_R_11 <= _GEN_57;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_12 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_12 <= _GEN_61;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_12 <= _GEN_61;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_12 <= 1'h0;
            end else begin
              in_live_in_valid_R_12 <= _GEN_61;
            end
          end else begin
            in_live_in_valid_R_12 <= _GEN_61;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_13 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_13 <= _GEN_65;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_13 <= _GEN_65;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_13 <= 1'h0;
            end else begin
              in_live_in_valid_R_13 <= _GEN_65;
            end
          end else begin
            in_live_in_valid_R_13 <= _GEN_65;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_14 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_14 <= _GEN_69;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_14 <= _GEN_69;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_14 <= 1'h0;
            end else begin
              in_live_in_valid_R_14 <= _GEN_69;
            end
          end else begin
            in_live_in_valid_R_14 <= _GEN_69;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_15 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_live_in_valid_R_15 <= _GEN_73;
      end else begin
        if (_T_115) begin
          in_live_in_valid_R_15 <= _GEN_73;
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_15 <= 1'h0;
            end else begin
              in_live_in_valid_R_15 <= _GEN_73;
            end
          end else begin
            in_live_in_valid_R_15 <= _GEN_73;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_66) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_66) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        in_carry_in_valid_R_0 <= _GEN_77;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_77;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_77;
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_77;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_77;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_0_0 <= _GEN_132;
        end else begin
          if (_T_70) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_0_0 <= _GEN_241;
          end else begin
            if (_T_70) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_70) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_1_0 <= _GEN_133;
        end else begin
          if (_T_71) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_1_0 <= _GEN_242;
          end else begin
            if (_T_71) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_71) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_2_0 <= _GEN_134;
        end else begin
          if (_T_72) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_2_0 <= _GEN_243;
          end else begin
            if (_T_72) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_72) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_3_0 <= _GEN_135;
        end else begin
          if (_T_73) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_3_0 <= _GEN_244;
          end else begin
            if (_T_73) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_73) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_4_0 <= _GEN_136;
        end else begin
          if (_T_74) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_4_0 <= _GEN_245;
          end else begin
            if (_T_74) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_74) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_5_0 <= _GEN_137;
        end else begin
          if (_T_75) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_5_0 <= _GEN_246;
          end else begin
            if (_T_75) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_75) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_6_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_6_0 <= _GEN_138;
        end else begin
          if (_T_76) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_6_0 <= _GEN_247;
          end else begin
            if (_T_76) begin
              out_live_in_valid_R_6_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_7_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_7_0 <= _GEN_139;
        end else begin
          if (_T_77) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_7_0 <= _GEN_248;
          end else begin
            if (_T_77) begin
              out_live_in_valid_R_7_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_77) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_8_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_8_0 <= _GEN_140;
        end else begin
          if (_T_78) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_8_0 <= _GEN_249;
          end else begin
            if (_T_78) begin
              out_live_in_valid_R_8_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_78) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_9_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_9_0 <= _GEN_141;
        end else begin
          if (_T_79) begin
            out_live_in_valid_R_9_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_9_0 <= _GEN_250;
          end else begin
            if (_T_79) begin
              out_live_in_valid_R_9_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_79) begin
            out_live_in_valid_R_9_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_10_0 <= _GEN_142;
        end else begin
          if (_T_80) begin
            out_live_in_valid_R_10_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_10_0 <= _GEN_251;
          end else begin
            if (_T_80) begin
              out_live_in_valid_R_10_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_80) begin
            out_live_in_valid_R_10_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_1 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_10_1 <= _GEN_143;
        end else begin
          if (_T_81) begin
            out_live_in_valid_R_10_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_10_1 <= _GEN_252;
          end else begin
            if (_T_81) begin
              out_live_in_valid_R_10_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_81) begin
            out_live_in_valid_R_10_1 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_2 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_10_2 <= _GEN_144;
        end else begin
          if (_T_82) begin
            out_live_in_valid_R_10_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_10_2 <= _GEN_253;
          end else begin
            if (_T_82) begin
              out_live_in_valid_R_10_2 <= 1'h0;
            end
          end
        end else begin
          if (_T_82) begin
            out_live_in_valid_R_10_2 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_3 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_10_3 <= _GEN_145;
        end else begin
          if (_T_83) begin
            out_live_in_valid_R_10_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_10_3 <= _GEN_254;
          end else begin
            if (_T_83) begin
              out_live_in_valid_R_10_3 <= 1'h0;
            end
          end
        end else begin
          if (_T_83) begin
            out_live_in_valid_R_10_3 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_4 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_10_4 <= _GEN_146;
        end else begin
          if (_T_84) begin
            out_live_in_valid_R_10_4 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_10_4 <= _GEN_255;
          end else begin
            if (_T_84) begin
              out_live_in_valid_R_10_4 <= 1'h0;
            end
          end
        end else begin
          if (_T_84) begin
            out_live_in_valid_R_10_4 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_5 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_10_5 <= _GEN_147;
        end else begin
          if (_T_85) begin
            out_live_in_valid_R_10_5 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_10_5 <= _GEN_256;
          end else begin
            if (_T_85) begin
              out_live_in_valid_R_10_5 <= 1'h0;
            end
          end
        end else begin
          if (_T_85) begin
            out_live_in_valid_R_10_5 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_6 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_10_6 <= _GEN_148;
        end else begin
          if (_T_86) begin
            out_live_in_valid_R_10_6 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_10_6 <= _GEN_257;
          end else begin
            if (_T_86) begin
              out_live_in_valid_R_10_6 <= 1'h0;
            end
          end
        end else begin
          if (_T_86) begin
            out_live_in_valid_R_10_6 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_7 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_10_7 <= _GEN_149;
        end else begin
          if (_T_87) begin
            out_live_in_valid_R_10_7 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_10_7 <= _GEN_258;
          end else begin
            if (_T_87) begin
              out_live_in_valid_R_10_7 <= 1'h0;
            end
          end
        end else begin
          if (_T_87) begin
            out_live_in_valid_R_10_7 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_8 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_10_8 <= _GEN_150;
        end else begin
          if (_T_88) begin
            out_live_in_valid_R_10_8 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_10_8 <= _GEN_259;
          end else begin
            if (_T_88) begin
              out_live_in_valid_R_10_8 <= 1'h0;
            end
          end
        end else begin
          if (_T_88) begin
            out_live_in_valid_R_10_8 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_11_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_11_0 <= _GEN_151;
        end else begin
          if (_T_89) begin
            out_live_in_valid_R_11_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_11_0 <= _GEN_260;
          end else begin
            if (_T_89) begin
              out_live_in_valid_R_11_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_89) begin
            out_live_in_valid_R_11_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_12_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_12_0 <= _GEN_152;
        end else begin
          if (_T_90) begin
            out_live_in_valid_R_12_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_12_0 <= _GEN_261;
          end else begin
            if (_T_90) begin
              out_live_in_valid_R_12_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_90) begin
            out_live_in_valid_R_12_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_13_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_13_0 <= _GEN_153;
        end else begin
          if (_T_91) begin
            out_live_in_valid_R_13_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_13_0 <= _GEN_262;
          end else begin
            if (_T_91) begin
              out_live_in_valid_R_13_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_91) begin
            out_live_in_valid_R_13_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_14_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_14_0 <= _GEN_154;
        end else begin
          if (_T_92) begin
            out_live_in_valid_R_14_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_14_0 <= _GEN_263;
          end else begin
            if (_T_92) begin
              out_live_in_valid_R_14_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_92) begin
            out_live_in_valid_R_14_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_15_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_live_in_valid_R_15_0 <= _GEN_155;
        end else begin
          if (_T_93) begin
            out_live_in_valid_R_15_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_live_in_valid_R_15_0 <= _GEN_264;
          end else begin
            if (_T_93) begin
              out_live_in_valid_R_15_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_93) begin
            out_live_in_valid_R_15_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_0_0 <= _GEN_83;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_0 <= _GEN_83;
            end
          end else begin
            out_live_in_fire_R_0_0 <= _GEN_83;
          end
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_83;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_1_0 <= _GEN_85;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_0 <= _GEN_85;
            end
          end else begin
            out_live_in_fire_R_1_0 <= _GEN_85;
          end
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_85;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_2_0 <= _GEN_87;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_2_0 <= _GEN_87;
            end
          end else begin
            out_live_in_fire_R_2_0 <= _GEN_87;
          end
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_87;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_3_0 <= _GEN_89;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_3_0 <= _GEN_89;
            end
          end else begin
            out_live_in_fire_R_3_0 <= _GEN_89;
          end
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_89;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_4_0 <= _GEN_91;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_4_0 <= _GEN_91;
            end
          end else begin
            out_live_in_fire_R_4_0 <= _GEN_91;
          end
        end else begin
          out_live_in_fire_R_4_0 <= _GEN_91;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_5_0 <= _GEN_93;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_5_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_5_0 <= _GEN_93;
            end
          end else begin
            out_live_in_fire_R_5_0 <= _GEN_93;
          end
        end else begin
          out_live_in_fire_R_5_0 <= _GEN_93;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_6_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_6_0 <= _GEN_95;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_6_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_6_0 <= _GEN_95;
            end
          end else begin
            out_live_in_fire_R_6_0 <= _GEN_95;
          end
        end else begin
          out_live_in_fire_R_6_0 <= _GEN_95;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_7_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_7_0 <= _GEN_97;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_7_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_7_0 <= _GEN_97;
            end
          end else begin
            out_live_in_fire_R_7_0 <= _GEN_97;
          end
        end else begin
          out_live_in_fire_R_7_0 <= _GEN_97;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_8_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_8_0 <= _GEN_99;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_8_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_8_0 <= _GEN_99;
            end
          end else begin
            out_live_in_fire_R_8_0 <= _GEN_99;
          end
        end else begin
          out_live_in_fire_R_8_0 <= _GEN_99;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_9_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_9_0 <= _GEN_101;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_9_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_9_0 <= _GEN_101;
            end
          end else begin
            out_live_in_fire_R_9_0 <= _GEN_101;
          end
        end else begin
          out_live_in_fire_R_9_0 <= _GEN_101;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_10_0 <= _GEN_103;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_0 <= _GEN_103;
            end
          end else begin
            out_live_in_fire_R_10_0 <= _GEN_103;
          end
        end else begin
          out_live_in_fire_R_10_0 <= _GEN_103;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_1 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_10_1 <= _GEN_105;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_1 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_1 <= _GEN_105;
            end
          end else begin
            out_live_in_fire_R_10_1 <= _GEN_105;
          end
        end else begin
          out_live_in_fire_R_10_1 <= _GEN_105;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_2 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_10_2 <= _GEN_107;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_2 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_2 <= _GEN_107;
            end
          end else begin
            out_live_in_fire_R_10_2 <= _GEN_107;
          end
        end else begin
          out_live_in_fire_R_10_2 <= _GEN_107;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_3 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_10_3 <= _GEN_109;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_3 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_3 <= _GEN_109;
            end
          end else begin
            out_live_in_fire_R_10_3 <= _GEN_109;
          end
        end else begin
          out_live_in_fire_R_10_3 <= _GEN_109;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_4 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_10_4 <= _GEN_111;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_4 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_4 <= _GEN_111;
            end
          end else begin
            out_live_in_fire_R_10_4 <= _GEN_111;
          end
        end else begin
          out_live_in_fire_R_10_4 <= _GEN_111;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_5 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_10_5 <= _GEN_113;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_5 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_5 <= _GEN_113;
            end
          end else begin
            out_live_in_fire_R_10_5 <= _GEN_113;
          end
        end else begin
          out_live_in_fire_R_10_5 <= _GEN_113;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_6 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_10_6 <= _GEN_115;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_6 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_6 <= _GEN_115;
            end
          end else begin
            out_live_in_fire_R_10_6 <= _GEN_115;
          end
        end else begin
          out_live_in_fire_R_10_6 <= _GEN_115;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_7 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_10_7 <= _GEN_117;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_7 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_7 <= _GEN_117;
            end
          end else begin
            out_live_in_fire_R_10_7 <= _GEN_117;
          end
        end else begin
          out_live_in_fire_R_10_7 <= _GEN_117;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_8 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_10_8 <= _GEN_119;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_8 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_8 <= _GEN_119;
            end
          end else begin
            out_live_in_fire_R_10_8 <= _GEN_119;
          end
        end else begin
          out_live_in_fire_R_10_8 <= _GEN_119;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_11_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_11_0 <= _GEN_121;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_11_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_11_0 <= _GEN_121;
            end
          end else begin
            out_live_in_fire_R_11_0 <= _GEN_121;
          end
        end else begin
          out_live_in_fire_R_11_0 <= _GEN_121;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_12_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_12_0 <= _GEN_123;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_12_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_12_0 <= _GEN_123;
            end
          end else begin
            out_live_in_fire_R_12_0 <= _GEN_123;
          end
        end else begin
          out_live_in_fire_R_12_0 <= _GEN_123;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_13_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_13_0 <= _GEN_125;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_13_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_13_0 <= _GEN_125;
            end
          end else begin
            out_live_in_fire_R_13_0 <= _GEN_125;
          end
        end else begin
          out_live_in_fire_R_13_0 <= _GEN_125;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_14_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_14_0 <= _GEN_127;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_14_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_14_0 <= _GEN_127;
            end
          end else begin
            out_live_in_fire_R_14_0 <= _GEN_127;
          end
        end else begin
          out_live_in_fire_R_14_0 <= _GEN_127;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_15_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        out_live_in_fire_R_15_0 <= _GEN_129;
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_15_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_15_0 <= _GEN_129;
            end
          end else begin
            out_live_in_fire_R_15_0 <= _GEN_129;
          end
        end else begin
          out_live_in_fire_R_15_0 <= _GEN_129;
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          out_carry_out_valid_R_0_0 <= _GEN_156;
        end else begin
          if (_T_94) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            out_carry_out_valid_R_0_0 <= _GEN_265;
          end else begin
            if (_T_94) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_94) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          active_loop_start_R_control <= _GEN_157;
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          active_loop_start_valid_R <= _GEN_159;
        end else begin
          if (_T_67) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            active_loop_start_valid_R <= _GEN_212;
          end else begin
            if (_T_67) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_67) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            active_loop_back_R_control <= _GEN_213;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          active_loop_back_valid_R <= _GEN_162;
        end else begin
          if (_T_68) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            active_loop_back_valid_R <= _GEN_215;
          end else begin
            if (_T_68) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_68) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 5'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          loop_exit_R_0_control <= _GEN_164;
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (!(loop_back_R_0_control)) begin
              loop_exit_R_0_control <= _GEN_207;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          if (enable_R_control) begin
            if (_T_69) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_69) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              if (_T_69) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              loop_exit_valid_R_0 <= _GEN_202;
            end
          end else begin
            if (_T_69) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_80;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_81;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_95) begin
        if (_T_111) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_115) begin
          if (_T_141) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_157) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_765 & _T_149) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOOP]   Loop_0: Restarted fired @ %d\n",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 932:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_771 & _T_149) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOOP]   Loop_0: Output fired @ %d ",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 950:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_771 & _T_149) begin
          $fwrite(32'h80000002,"\n"); // @[LoopBlock.scala 955:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LoopBlockNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_InLiveIn_0_ready,
  input         io_InLiveIn_0_valid,
  input  [31:0] io_InLiveIn_0_bits_data,
  output        io_InLiveIn_1_ready,
  input         io_InLiveIn_1_valid,
  input  [31:0] io_InLiveIn_1_bits_data,
  output        io_InLiveIn_2_ready,
  input         io_InLiveIn_2_valid,
  input  [4:0]  io_InLiveIn_2_bits_taskID,
  input  [31:0] io_InLiveIn_2_bits_data,
  output        io_InLiveIn_3_ready,
  input         io_InLiveIn_3_valid,
  input         io_InLiveIn_3_bits_predicate,
  input  [4:0]  io_InLiveIn_3_bits_taskID,
  input  [31:0] io_InLiveIn_3_bits_data,
  output        io_InLiveIn_4_ready,
  input         io_InLiveIn_4_valid,
  input  [4:0]  io_InLiveIn_4_bits_taskID,
  input  [31:0] io_InLiveIn_4_bits_data,
  output        io_InLiveIn_5_ready,
  input         io_InLiveIn_5_valid,
  input         io_InLiveIn_5_bits_predicate,
  input  [4:0]  io_InLiveIn_5_bits_taskID,
  input  [31:0] io_InLiveIn_5_bits_data,
  output        io_InLiveIn_6_ready,
  input         io_InLiveIn_6_valid,
  input         io_InLiveIn_6_bits_predicate,
  input  [4:0]  io_InLiveIn_6_bits_taskID,
  input  [31:0] io_InLiveIn_6_bits_data,
  output        io_InLiveIn_7_ready,
  input         io_InLiveIn_7_valid,
  input         io_InLiveIn_7_bits_predicate,
  input  [4:0]  io_InLiveIn_7_bits_taskID,
  input  [31:0] io_InLiveIn_7_bits_data,
  output        io_InLiveIn_8_ready,
  input         io_InLiveIn_8_valid,
  input         io_InLiveIn_8_bits_predicate,
  input  [4:0]  io_InLiveIn_8_bits_taskID,
  input  [31:0] io_InLiveIn_8_bits_data,
  output        io_InLiveIn_9_ready,
  input         io_InLiveIn_9_valid,
  input         io_InLiveIn_9_bits_predicate,
  input  [4:0]  io_InLiveIn_9_bits_taskID,
  input  [31:0] io_InLiveIn_9_bits_data,
  output        io_InLiveIn_10_ready,
  input         io_InLiveIn_10_valid,
  input         io_InLiveIn_10_bits_predicate,
  input  [4:0]  io_InLiveIn_10_bits_taskID,
  input  [31:0] io_InLiveIn_10_bits_data,
  output        io_InLiveIn_11_ready,
  input         io_InLiveIn_11_valid,
  input         io_InLiveIn_11_bits_predicate,
  input  [4:0]  io_InLiveIn_11_bits_taskID,
  input  [31:0] io_InLiveIn_11_bits_data,
  output        io_InLiveIn_12_ready,
  input         io_InLiveIn_12_valid,
  input         io_InLiveIn_12_bits_predicate,
  input  [4:0]  io_InLiveIn_12_bits_taskID,
  input  [31:0] io_InLiveIn_12_bits_data,
  input         io_OutLiveIn_field12_0_ready,
  output        io_OutLiveIn_field12_0_valid,
  output        io_OutLiveIn_field12_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field12_0_bits_taskID,
  output [31:0] io_OutLiveIn_field12_0_bits_data,
  input         io_OutLiveIn_field11_0_ready,
  output        io_OutLiveIn_field11_0_valid,
  output        io_OutLiveIn_field11_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field11_0_bits_taskID,
  output [31:0] io_OutLiveIn_field11_0_bits_data,
  input         io_OutLiveIn_field10_0_ready,
  output        io_OutLiveIn_field10_0_valid,
  output        io_OutLiveIn_field10_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field10_0_bits_taskID,
  output [31:0] io_OutLiveIn_field10_0_bits_data,
  input         io_OutLiveIn_field9_0_ready,
  output        io_OutLiveIn_field9_0_valid,
  output        io_OutLiveIn_field9_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field9_0_bits_taskID,
  output [31:0] io_OutLiveIn_field9_0_bits_data,
  input         io_OutLiveIn_field8_0_ready,
  output        io_OutLiveIn_field8_0_valid,
  output        io_OutLiveIn_field8_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field8_0_bits_taskID,
  output [31:0] io_OutLiveIn_field8_0_bits_data,
  input         io_OutLiveIn_field7_0_ready,
  output        io_OutLiveIn_field7_0_valid,
  output        io_OutLiveIn_field7_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field7_0_bits_taskID,
  output [31:0] io_OutLiveIn_field7_0_bits_data,
  input         io_OutLiveIn_field6_0_ready,
  output        io_OutLiveIn_field6_0_valid,
  output        io_OutLiveIn_field6_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field6_0_bits_taskID,
  output [31:0] io_OutLiveIn_field6_0_bits_data,
  input         io_OutLiveIn_field5_0_ready,
  output        io_OutLiveIn_field5_0_valid,
  output        io_OutLiveIn_field5_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field5_0_bits_taskID,
  output [31:0] io_OutLiveIn_field5_0_bits_data,
  input         io_OutLiveIn_field4_0_ready,
  output        io_OutLiveIn_field4_0_valid,
  output [4:0]  io_OutLiveIn_field4_0_bits_taskID,
  output [31:0] io_OutLiveIn_field4_0_bits_data,
  input         io_OutLiveIn_field3_0_ready,
  output        io_OutLiveIn_field3_0_valid,
  output        io_OutLiveIn_field3_0_bits_predicate,
  output [4:0]  io_OutLiveIn_field3_0_bits_taskID,
  output [31:0] io_OutLiveIn_field3_0_bits_data,
  input         io_OutLiveIn_field2_0_ready,
  output        io_OutLiveIn_field2_0_valid,
  output [4:0]  io_OutLiveIn_field2_0_bits_taskID,
  output [31:0] io_OutLiveIn_field2_0_bits_data,
  input         io_OutLiveIn_field1_0_ready,
  output        io_OutLiveIn_field1_0_valid,
  output [31:0] io_OutLiveIn_field1_0_bits_data,
  input         io_OutLiveIn_field1_1_ready,
  output        io_OutLiveIn_field1_1_valid,
  output [31:0] io_OutLiveIn_field1_1_bits_data,
  input         io_OutLiveIn_field1_2_ready,
  output        io_OutLiveIn_field1_2_valid,
  output [31:0] io_OutLiveIn_field1_2_bits_data,
  input         io_OutLiveIn_field0_0_ready,
  output        io_OutLiveIn_field0_0_valid,
  output [31:0] io_OutLiveIn_field0_0_bits_data,
  input         io_OutLiveIn_field0_1_ready,
  output        io_OutLiveIn_field0_1_valid,
  output [31:0] io_OutLiveIn_field0_1_bits_data,
  input         io_OutLiveIn_field0_2_ready,
  output        io_OutLiveIn_field0_2_valid,
  output [31:0] io_OutLiveIn_field0_2_bits_data,
  input         io_activate_loop_start_ready,
  output        io_activate_loop_start_valid,
  output [4:0]  io_activate_loop_start_bits_taskID,
  output        io_activate_loop_start_bits_control,
  input         io_activate_loop_back_ready,
  output        io_activate_loop_back_valid,
  output [4:0]  io_activate_loop_back_bits_taskID,
  output        io_activate_loop_back_bits_control,
  output        io_loopBack_0_ready,
  input         io_loopBack_0_valid,
  input  [4:0]  io_loopBack_0_bits_taskID,
  input         io_loopBack_0_bits_control,
  output        io_loopFinish_0_ready,
  input         io_loopFinish_0_valid,
  input         io_loopFinish_0_bits_control,
  output        io_CarryDepenIn_0_ready,
  input         io_CarryDepenIn_0_valid,
  input  [4:0]  io_CarryDepenIn_0_bits_taskID,
  input  [31:0] io_CarryDepenIn_0_bits_data,
  input         io_CarryDepenOut_field0_0_ready,
  output        io_CarryDepenOut_field0_0_valid,
  output [4:0]  io_CarryDepenOut_field0_0_bits_taskID,
  output [31:0] io_CarryDepenOut_field0_0_bits_data,
  input         io_loopExit_0_ready,
  output        io_loopExit_0_valid,
  output [4:0]  io_loopExit_0_bits_taskID,
  output        io_loopExit_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_1;
  reg  enable_R_control; // @[LoopBlock.scala 528:25]
  reg [31:0] _RAND_2;
  reg  enable_valid_R; // @[LoopBlock.scala 529:31]
  reg [31:0] _RAND_3;
  reg [4:0] loop_back_R_0_taskID; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_4;
  reg  loop_back_R_0_control; // @[LoopBlock.scala 531:50]
  reg [31:0] _RAND_5;
  reg  loop_back_valid_R_0; // @[LoopBlock.scala 532:56]
  reg [31:0] _RAND_6;
  reg  loop_finish_R_0_control; // @[LoopBlock.scala 534:54]
  reg [31:0] _RAND_7;
  reg  loop_finish_valid_R_0; // @[LoopBlock.scala 535:60]
  reg [31:0] _RAND_8;
  reg [31:0] in_live_in_R_0_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_9;
  reg [31:0] in_live_in_R_1_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_10;
  reg [4:0] in_live_in_R_2_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_11;
  reg [31:0] in_live_in_R_2_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_12;
  reg  in_live_in_R_3_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_13;
  reg [4:0] in_live_in_R_3_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_14;
  reg [31:0] in_live_in_R_3_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_15;
  reg [4:0] in_live_in_R_4_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_16;
  reg [31:0] in_live_in_R_4_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_17;
  reg  in_live_in_R_5_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_18;
  reg [4:0] in_live_in_R_5_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_19;
  reg [31:0] in_live_in_R_5_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_20;
  reg  in_live_in_R_6_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_21;
  reg [4:0] in_live_in_R_6_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_22;
  reg [31:0] in_live_in_R_6_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_23;
  reg  in_live_in_R_7_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_24;
  reg [4:0] in_live_in_R_7_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_25;
  reg [31:0] in_live_in_R_7_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_26;
  reg  in_live_in_R_8_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_27;
  reg [4:0] in_live_in_R_8_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_28;
  reg [31:0] in_live_in_R_8_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_29;
  reg  in_live_in_R_9_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_30;
  reg [4:0] in_live_in_R_9_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_31;
  reg [31:0] in_live_in_R_9_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_32;
  reg  in_live_in_R_10_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_33;
  reg [4:0] in_live_in_R_10_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_34;
  reg [31:0] in_live_in_R_10_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_35;
  reg  in_live_in_R_11_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_36;
  reg [4:0] in_live_in_R_11_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_37;
  reg [31:0] in_live_in_R_11_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_38;
  reg  in_live_in_R_12_predicate; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_39;
  reg [4:0] in_live_in_R_12_taskID; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_40;
  reg [31:0] in_live_in_R_12_data; // @[LoopBlock.scala 537:53]
  reg [31:0] _RAND_41;
  reg  in_live_in_valid_R_0; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_42;
  reg  in_live_in_valid_R_1; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_43;
  reg  in_live_in_valid_R_2; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_44;
  reg  in_live_in_valid_R_3; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_45;
  reg  in_live_in_valid_R_4; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_46;
  reg  in_live_in_valid_R_5; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_47;
  reg  in_live_in_valid_R_6; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_48;
  reg  in_live_in_valid_R_7; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_49;
  reg  in_live_in_valid_R_8; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_50;
  reg  in_live_in_valid_R_9; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_51;
  reg  in_live_in_valid_R_10; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_52;
  reg  in_live_in_valid_R_11; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_53;
  reg  in_live_in_valid_R_12; // @[LoopBlock.scala 538:59]
  reg [31:0] _RAND_54;
  reg [4:0] in_carry_in_R_0_taskID; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_55;
  reg [31:0] in_carry_in_R_0_data; // @[LoopBlock.scala 540:56]
  reg [31:0] _RAND_56;
  reg  in_carry_in_valid_R_0; // @[LoopBlock.scala 541:62]
  reg [31:0] _RAND_57;
  reg  out_live_in_valid_R_0_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_58;
  reg  out_live_in_valid_R_0_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_59;
  reg  out_live_in_valid_R_0_2; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_60;
  reg  out_live_in_valid_R_1_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_61;
  reg  out_live_in_valid_R_1_1; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_62;
  reg  out_live_in_valid_R_1_2; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_63;
  reg  out_live_in_valid_R_2_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_64;
  reg  out_live_in_valid_R_3_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_65;
  reg  out_live_in_valid_R_4_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_66;
  reg  out_live_in_valid_R_5_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_67;
  reg  out_live_in_valid_R_6_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_68;
  reg  out_live_in_valid_R_7_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_69;
  reg  out_live_in_valid_R_8_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_70;
  reg  out_live_in_valid_R_9_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_71;
  reg  out_live_in_valid_R_10_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_72;
  reg  out_live_in_valid_R_11_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_73;
  reg  out_live_in_valid_R_12_0; // @[LoopBlock.scala 553:47]
  reg [31:0] _RAND_74;
  reg  out_live_in_fire_R_0_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_75;
  reg  out_live_in_fire_R_0_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_76;
  reg  out_live_in_fire_R_0_2; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_77;
  reg  out_live_in_fire_R_1_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_78;
  reg  out_live_in_fire_R_1_1; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_79;
  reg  out_live_in_fire_R_1_2; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_80;
  reg  out_live_in_fire_R_2_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_81;
  reg  out_live_in_fire_R_3_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_82;
  reg  out_live_in_fire_R_4_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_83;
  reg  out_live_in_fire_R_5_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_84;
  reg  out_live_in_fire_R_6_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_85;
  reg  out_live_in_fire_R_7_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_86;
  reg  out_live_in_fire_R_8_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_87;
  reg  out_live_in_fire_R_9_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_88;
  reg  out_live_in_fire_R_10_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_89;
  reg  out_live_in_fire_R_11_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_90;
  reg  out_live_in_fire_R_12_0; // @[LoopBlock.scala 557:47]
  reg [31:0] _RAND_91;
  reg  out_carry_out_valid_R_0_0; // @[LoopBlock.scala 573:44]
  reg [31:0] _RAND_92;
  reg [4:0] active_loop_start_R_taskID; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_93;
  reg  active_loop_start_R_control; // @[LoopBlock.scala 581:36]
  reg [31:0] _RAND_94;
  reg  active_loop_start_valid_R; // @[LoopBlock.scala 582:42]
  reg [31:0] _RAND_95;
  reg [4:0] active_loop_back_R_taskID; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_96;
  reg  active_loop_back_R_control; // @[LoopBlock.scala 584:35]
  reg [31:0] _RAND_97;
  reg  active_loop_back_valid_R; // @[LoopBlock.scala 585:41]
  reg [31:0] _RAND_98;
  reg [4:0] loop_exit_R_0_taskID; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_99;
  reg  loop_exit_R_0_control; // @[LoopBlock.scala 587:47]
  reg [31:0] _RAND_100;
  reg  loop_exit_valid_R_0; // @[LoopBlock.scala 588:53]
  reg [31:0] _RAND_101;
  reg  loop_exit_fire_R_0; // @[LoopBlock.scala 589:52]
  reg [31:0] _RAND_102;
  wire  _T_25; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[LoopBlock.scala 596:26]
  wire  _T_27; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[LoopBlock.scala 603:33]
  wire [4:0] _GEN_5; // @[LoopBlock.scala 603:33]
  wire  _GEN_6; // @[LoopBlock.scala 603:33]
  wire  _T_29; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[LoopBlock.scala 612:35]
  wire  _GEN_9; // @[LoopBlock.scala 612:35]
  wire  _T_31; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[LoopBlock.scala 623:33]
  wire  _T_33; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[LoopBlock.scala 623:33]
  wire  _T_35; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[LoopBlock.scala 623:33]
  wire  _T_37; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[LoopBlock.scala 623:33]
  wire  _T_39; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[LoopBlock.scala 623:33]
  wire  _T_41; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[LoopBlock.scala 623:33]
  wire  _T_43; // @[Decoupled.scala 40:37]
  wire  _GEN_37; // @[LoopBlock.scala 623:33]
  wire  _T_45; // @[Decoupled.scala 40:37]
  wire  _GEN_41; // @[LoopBlock.scala 623:33]
  wire  _T_47; // @[Decoupled.scala 40:37]
  wire  _GEN_45; // @[LoopBlock.scala 623:33]
  wire  _T_49; // @[Decoupled.scala 40:37]
  wire  _GEN_49; // @[LoopBlock.scala 623:33]
  wire  _T_51; // @[Decoupled.scala 40:37]
  wire  _GEN_53; // @[LoopBlock.scala 623:33]
  wire  _T_53; // @[Decoupled.scala 40:37]
  wire  _GEN_57; // @[LoopBlock.scala 623:33]
  wire  _T_55; // @[Decoupled.scala 40:37]
  wire  _GEN_61; // @[LoopBlock.scala 623:33]
  wire  _T_57; // @[Decoupled.scala 40:37]
  wire  _GEN_65; // @[LoopBlock.scala 641:37]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire  _GEN_66; // @[LoopBlock.scala 704:39]
  wire  _T_59; // @[Decoupled.scala 40:37]
  wire  _GEN_67; // @[LoopBlock.scala 708:38]
  wire  _T_60; // @[Decoupled.scala 40:37]
  wire  _GEN_68; // @[LoopBlock.scala 713:33]
  wire  _GEN_69; // @[LoopBlock.scala 713:33]
  wire  _T_61; // @[Decoupled.scala 40:37]
  wire  _GEN_70; // @[LoopBlock.scala 722:57]
  wire  _GEN_71; // @[LoopBlock.scala 722:57]
  wire  _T_62; // @[Decoupled.scala 40:37]
  wire  _GEN_72; // @[LoopBlock.scala 722:57]
  wire  _GEN_73; // @[LoopBlock.scala 722:57]
  wire  _T_63; // @[Decoupled.scala 40:37]
  wire  _GEN_74; // @[LoopBlock.scala 722:57]
  wire  _GEN_75; // @[LoopBlock.scala 722:57]
  wire  _T_64; // @[Decoupled.scala 40:37]
  wire  _GEN_76; // @[LoopBlock.scala 722:57]
  wire  _GEN_77; // @[LoopBlock.scala 722:57]
  wire  _T_65; // @[Decoupled.scala 40:37]
  wire  _GEN_78; // @[LoopBlock.scala 722:57]
  wire  _GEN_79; // @[LoopBlock.scala 722:57]
  wire  _T_66; // @[Decoupled.scala 40:37]
  wire  _GEN_80; // @[LoopBlock.scala 722:57]
  wire  _GEN_81; // @[LoopBlock.scala 722:57]
  wire  _T_67; // @[Decoupled.scala 40:37]
  wire  _GEN_82; // @[LoopBlock.scala 722:57]
  wire  _GEN_83; // @[LoopBlock.scala 722:57]
  wire  _T_68; // @[Decoupled.scala 40:37]
  wire  _GEN_84; // @[LoopBlock.scala 722:57]
  wire  _GEN_85; // @[LoopBlock.scala 722:57]
  wire  _T_69; // @[Decoupled.scala 40:37]
  wire  _GEN_86; // @[LoopBlock.scala 722:57]
  wire  _GEN_87; // @[LoopBlock.scala 722:57]
  wire  _T_70; // @[Decoupled.scala 40:37]
  wire  _GEN_88; // @[LoopBlock.scala 722:57]
  wire  _GEN_89; // @[LoopBlock.scala 722:57]
  wire  _T_71; // @[Decoupled.scala 40:37]
  wire  _GEN_90; // @[LoopBlock.scala 722:57]
  wire  _GEN_91; // @[LoopBlock.scala 722:57]
  wire  _T_72; // @[Decoupled.scala 40:37]
  wire  _GEN_92; // @[LoopBlock.scala 722:57]
  wire  _GEN_93; // @[LoopBlock.scala 722:57]
  wire  _T_73; // @[Decoupled.scala 40:37]
  wire  _GEN_94; // @[LoopBlock.scala 722:57]
  wire  _GEN_95; // @[LoopBlock.scala 722:57]
  wire  _T_74; // @[Decoupled.scala 40:37]
  wire  _GEN_96; // @[LoopBlock.scala 722:57]
  wire  _GEN_97; // @[LoopBlock.scala 722:57]
  wire  _T_75; // @[Decoupled.scala 40:37]
  wire  _GEN_98; // @[LoopBlock.scala 722:57]
  wire  _GEN_99; // @[LoopBlock.scala 722:57]
  wire  _T_76; // @[Decoupled.scala 40:37]
  wire  _GEN_100; // @[LoopBlock.scala 722:57]
  wire  _GEN_101; // @[LoopBlock.scala 722:57]
  wire  _T_77; // @[Decoupled.scala 40:37]
  wire  _GEN_102; // @[LoopBlock.scala 722:57]
  wire  _GEN_103; // @[LoopBlock.scala 722:57]
  wire  _T_78; // @[Decoupled.scala 40:37]
  wire  _GEN_104; // @[LoopBlock.scala 742:61]
  reg [1:0] state; // @[LoopBlock.scala 861:22]
  reg [31:0] _RAND_103;
  wire  _T_79; // @[Conditional.scala 37:30]
  wire  _T_80; // @[LoopBlock.scala 765:35]
  wire  _T_81; // @[LoopBlock.scala 765:35]
  wire  _T_82; // @[LoopBlock.scala 765:35]
  wire  _T_83; // @[LoopBlock.scala 765:35]
  wire  _T_84; // @[LoopBlock.scala 765:35]
  wire  _T_85; // @[LoopBlock.scala 765:35]
  wire  _T_86; // @[LoopBlock.scala 765:35]
  wire  _T_87; // @[LoopBlock.scala 765:35]
  wire  _T_88; // @[LoopBlock.scala 765:35]
  wire  _T_89; // @[LoopBlock.scala 765:35]
  wire  _T_90; // @[LoopBlock.scala 765:35]
  wire  _T_91; // @[LoopBlock.scala 765:35]
  wire  _T_92; // @[LoopBlock.scala 869:28]
  wire  _GEN_106; // @[LoopBlock.scala 870:26]
  wire  _GEN_107; // @[LoopBlock.scala 870:26]
  wire  _GEN_108; // @[LoopBlock.scala 870:26]
  wire  _GEN_109; // @[LoopBlock.scala 870:26]
  wire  _GEN_110; // @[LoopBlock.scala 870:26]
  wire  _GEN_111; // @[LoopBlock.scala 870:26]
  wire  _GEN_112; // @[LoopBlock.scala 870:26]
  wire  _GEN_113; // @[LoopBlock.scala 870:26]
  wire  _GEN_114; // @[LoopBlock.scala 870:26]
  wire  _GEN_115; // @[LoopBlock.scala 870:26]
  wire  _GEN_116; // @[LoopBlock.scala 870:26]
  wire  _GEN_117; // @[LoopBlock.scala 870:26]
  wire  _GEN_118; // @[LoopBlock.scala 870:26]
  wire  _GEN_119; // @[LoopBlock.scala 870:26]
  wire  _GEN_120; // @[LoopBlock.scala 870:26]
  wire  _GEN_121; // @[LoopBlock.scala 870:26]
  wire  _GEN_122; // @[LoopBlock.scala 870:26]
  wire  _GEN_123; // @[LoopBlock.scala 870:26]
  wire  _GEN_124; // @[LoopBlock.scala 870:26]
  wire  _GEN_126; // @[LoopBlock.scala 870:26]
  wire  _GEN_129; // @[LoopBlock.scala 870:26]
  wire  _GEN_131; // @[LoopBlock.scala 870:26]
  wire  _T_96; // @[Conditional.scala 37:30]
  wire  _T_97; // @[LoopBlock.scala 898:30]
  wire  _T_99; // @[LoopBlock.scala 825:65]
  wire  _T_100; // @[LoopBlock.scala 825:65]
  wire  _T_101; // @[LoopBlock.scala 825:65]
  wire  _T_102; // @[LoopBlock.scala 825:65]
  wire  _T_103; // @[LoopBlock.scala 828:26]
  wire  _T_104; // @[LoopBlock.scala 828:26]
  wire  _T_105; // @[LoopBlock.scala 828:26]
  wire  _T_106; // @[LoopBlock.scala 828:26]
  wire  _T_107; // @[LoopBlock.scala 828:26]
  wire  _T_108; // @[LoopBlock.scala 828:26]
  wire  _T_109; // @[LoopBlock.scala 828:26]
  wire  _T_110; // @[LoopBlock.scala 828:26]
  wire  _T_111; // @[LoopBlock.scala 828:26]
  wire  _T_112; // @[LoopBlock.scala 828:26]
  wire  _T_113; // @[LoopBlock.scala 828:26]
  wire  _T_114; // @[LoopBlock.scala 828:26]
  wire  _T_115; // @[LoopBlock.scala 899:29]
  wire  _T_122; // @[LoopBlock.scala 932:19]
  wire  _T_123; // @[LoopBlock.scala 932:19]
  wire  _GEN_162; // @[LoopBlock.scala 936:64]
  wire  _GEN_165; // @[LoopBlock.scala 936:64]
  wire  _GEN_167; // @[LoopBlock.scala 936:64]
  wire  _GEN_172; // @[LoopBlock.scala 903:56]
  wire  _GEN_173; // @[LoopBlock.scala 903:56]
  wire  _GEN_175; // @[LoopBlock.scala 903:56]
  wire  _GEN_194; // @[LoopBlock.scala 903:56]
  wire  _GEN_195; // @[LoopBlock.scala 903:56]
  wire  _GEN_196; // @[LoopBlock.scala 903:56]
  wire  _GEN_197; // @[LoopBlock.scala 903:56]
  wire  _GEN_198; // @[LoopBlock.scala 903:56]
  wire  _GEN_199; // @[LoopBlock.scala 903:56]
  wire  _GEN_200; // @[LoopBlock.scala 903:56]
  wire  _GEN_201; // @[LoopBlock.scala 903:56]
  wire  _GEN_202; // @[LoopBlock.scala 903:56]
  wire  _GEN_203; // @[LoopBlock.scala 903:56]
  wire  _GEN_204; // @[LoopBlock.scala 903:56]
  wire  _GEN_205; // @[LoopBlock.scala 903:56]
  wire  _GEN_206; // @[LoopBlock.scala 903:56]
  wire  _GEN_207; // @[LoopBlock.scala 903:56]
  wire  _GEN_208; // @[LoopBlock.scala 903:56]
  wire  _GEN_209; // @[LoopBlock.scala 903:56]
  wire  _GEN_210; // @[LoopBlock.scala 903:56]
  wire  _GEN_211; // @[LoopBlock.scala 903:56]
  wire  _T_131; // @[Conditional.scala 37:30]
  wire  _GEN_618; // @[LoopBlock.scala 932:19]
  wire  _GEN_619; // @[LoopBlock.scala 932:19]
  wire  _GEN_620; // @[LoopBlock.scala 932:19]
  wire  _GEN_621; // @[LoopBlock.scala 932:19]
  wire  _GEN_625; // @[LoopBlock.scala 950:19]
  wire  _GEN_626; // @[LoopBlock.scala 950:19]
  wire  _GEN_627; // @[LoopBlock.scala 950:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_25 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_25 | enable_valid_R; // @[LoopBlock.scala 596:26]
  assign _T_27 = io_loopBack_0_ready & io_loopBack_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_27 ? io_loopBack_0_bits_control : loop_back_R_0_control; // @[LoopBlock.scala 603:33]
  assign _GEN_5 = _T_27 ? io_loopBack_0_bits_taskID : loop_back_R_0_taskID; // @[LoopBlock.scala 603:33]
  assign _GEN_6 = _T_27 | loop_back_valid_R_0; // @[LoopBlock.scala 603:33]
  assign _T_29 = io_loopFinish_0_ready & io_loopFinish_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_29 ? io_loopFinish_0_bits_control : loop_finish_R_0_control; // @[LoopBlock.scala 612:35]
  assign _GEN_9 = _T_29 | loop_finish_valid_R_0; // @[LoopBlock.scala 612:35]
  assign _T_31 = io_InLiveIn_0_ready & io_InLiveIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_31 | in_live_in_valid_R_0; // @[LoopBlock.scala 623:33]
  assign _T_33 = io_InLiveIn_1_ready & io_InLiveIn_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_33 | in_live_in_valid_R_1; // @[LoopBlock.scala 623:33]
  assign _T_35 = io_InLiveIn_2_ready & io_InLiveIn_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_35 | in_live_in_valid_R_2; // @[LoopBlock.scala 623:33]
  assign _T_37 = io_InLiveIn_3_ready & io_InLiveIn_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_37 | in_live_in_valid_R_3; // @[LoopBlock.scala 623:33]
  assign _T_39 = io_InLiveIn_4_ready & io_InLiveIn_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_39 | in_live_in_valid_R_4; // @[LoopBlock.scala 623:33]
  assign _T_41 = io_InLiveIn_5_ready & io_InLiveIn_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_41 | in_live_in_valid_R_5; // @[LoopBlock.scala 623:33]
  assign _T_43 = io_InLiveIn_6_ready & io_InLiveIn_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_37 = _T_43 | in_live_in_valid_R_6; // @[LoopBlock.scala 623:33]
  assign _T_45 = io_InLiveIn_7_ready & io_InLiveIn_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_41 = _T_45 | in_live_in_valid_R_7; // @[LoopBlock.scala 623:33]
  assign _T_47 = io_InLiveIn_8_ready & io_InLiveIn_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_45 = _T_47 | in_live_in_valid_R_8; // @[LoopBlock.scala 623:33]
  assign _T_49 = io_InLiveIn_9_ready & io_InLiveIn_9_valid; // @[Decoupled.scala 40:37]
  assign _GEN_49 = _T_49 | in_live_in_valid_R_9; // @[LoopBlock.scala 623:33]
  assign _T_51 = io_InLiveIn_10_ready & io_InLiveIn_10_valid; // @[Decoupled.scala 40:37]
  assign _GEN_53 = _T_51 | in_live_in_valid_R_10; // @[LoopBlock.scala 623:33]
  assign _T_53 = io_InLiveIn_11_ready & io_InLiveIn_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_57 = _T_53 | in_live_in_valid_R_11; // @[LoopBlock.scala 623:33]
  assign _T_55 = io_InLiveIn_12_ready & io_InLiveIn_12_valid; // @[Decoupled.scala 40:37]
  assign _GEN_61 = _T_55 | in_live_in_valid_R_12; // @[LoopBlock.scala 623:33]
  assign _T_57 = io_CarryDepenIn_0_ready & io_CarryDepenIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_65 = _T_57 | in_carry_in_valid_R_0; // @[LoopBlock.scala 641:37]
  assign _T_58 = io_activate_loop_start_ready & io_activate_loop_start_valid; // @[Decoupled.scala 40:37]
  assign _GEN_66 = _T_58 ? 1'h0 : active_loop_start_valid_R; // @[LoopBlock.scala 704:39]
  assign _T_59 = io_activate_loop_back_ready & io_activate_loop_back_valid; // @[Decoupled.scala 40:37]
  assign _GEN_67 = _T_59 ? 1'h0 : active_loop_back_valid_R; // @[LoopBlock.scala 708:38]
  assign _T_60 = io_loopExit_0_ready & io_loopExit_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_68 = _T_60 ? 1'h0 : loop_exit_valid_R_0; // @[LoopBlock.scala 713:33]
  assign _GEN_69 = _T_60 | loop_exit_fire_R_0; // @[LoopBlock.scala 713:33]
  assign _T_61 = io_OutLiveIn_field0_0_ready & io_OutLiveIn_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_70 = _T_61 ? 1'h0 : out_live_in_valid_R_0_0; // @[LoopBlock.scala 722:57]
  assign _GEN_71 = _T_61 | out_live_in_fire_R_0_0; // @[LoopBlock.scala 722:57]
  assign _T_62 = io_OutLiveIn_field0_1_ready & io_OutLiveIn_field0_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_72 = _T_62 ? 1'h0 : out_live_in_valid_R_0_1; // @[LoopBlock.scala 722:57]
  assign _GEN_73 = _T_62 | out_live_in_fire_R_0_1; // @[LoopBlock.scala 722:57]
  assign _T_63 = io_OutLiveIn_field0_2_ready & io_OutLiveIn_field0_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_74 = _T_63 ? 1'h0 : out_live_in_valid_R_0_2; // @[LoopBlock.scala 722:57]
  assign _GEN_75 = _T_63 | out_live_in_fire_R_0_2; // @[LoopBlock.scala 722:57]
  assign _T_64 = io_OutLiveIn_field1_0_ready & io_OutLiveIn_field1_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_76 = _T_64 ? 1'h0 : out_live_in_valid_R_1_0; // @[LoopBlock.scala 722:57]
  assign _GEN_77 = _T_64 | out_live_in_fire_R_1_0; // @[LoopBlock.scala 722:57]
  assign _T_65 = io_OutLiveIn_field1_1_ready & io_OutLiveIn_field1_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_78 = _T_65 ? 1'h0 : out_live_in_valid_R_1_1; // @[LoopBlock.scala 722:57]
  assign _GEN_79 = _T_65 | out_live_in_fire_R_1_1; // @[LoopBlock.scala 722:57]
  assign _T_66 = io_OutLiveIn_field1_2_ready & io_OutLiveIn_field1_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_80 = _T_66 ? 1'h0 : out_live_in_valid_R_1_2; // @[LoopBlock.scala 722:57]
  assign _GEN_81 = _T_66 | out_live_in_fire_R_1_2; // @[LoopBlock.scala 722:57]
  assign _T_67 = io_OutLiveIn_field2_0_ready & io_OutLiveIn_field2_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_82 = _T_67 ? 1'h0 : out_live_in_valid_R_2_0; // @[LoopBlock.scala 722:57]
  assign _GEN_83 = _T_67 | out_live_in_fire_R_2_0; // @[LoopBlock.scala 722:57]
  assign _T_68 = io_OutLiveIn_field3_0_ready & io_OutLiveIn_field3_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_84 = _T_68 ? 1'h0 : out_live_in_valid_R_3_0; // @[LoopBlock.scala 722:57]
  assign _GEN_85 = _T_68 | out_live_in_fire_R_3_0; // @[LoopBlock.scala 722:57]
  assign _T_69 = io_OutLiveIn_field4_0_ready & io_OutLiveIn_field4_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_86 = _T_69 ? 1'h0 : out_live_in_valid_R_4_0; // @[LoopBlock.scala 722:57]
  assign _GEN_87 = _T_69 | out_live_in_fire_R_4_0; // @[LoopBlock.scala 722:57]
  assign _T_70 = io_OutLiveIn_field5_0_ready & io_OutLiveIn_field5_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_88 = _T_70 ? 1'h0 : out_live_in_valid_R_5_0; // @[LoopBlock.scala 722:57]
  assign _GEN_89 = _T_70 | out_live_in_fire_R_5_0; // @[LoopBlock.scala 722:57]
  assign _T_71 = io_OutLiveIn_field6_0_ready & io_OutLiveIn_field6_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_90 = _T_71 ? 1'h0 : out_live_in_valid_R_6_0; // @[LoopBlock.scala 722:57]
  assign _GEN_91 = _T_71 | out_live_in_fire_R_6_0; // @[LoopBlock.scala 722:57]
  assign _T_72 = io_OutLiveIn_field7_0_ready & io_OutLiveIn_field7_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_92 = _T_72 ? 1'h0 : out_live_in_valid_R_7_0; // @[LoopBlock.scala 722:57]
  assign _GEN_93 = _T_72 | out_live_in_fire_R_7_0; // @[LoopBlock.scala 722:57]
  assign _T_73 = io_OutLiveIn_field8_0_ready & io_OutLiveIn_field8_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_94 = _T_73 ? 1'h0 : out_live_in_valid_R_8_0; // @[LoopBlock.scala 722:57]
  assign _GEN_95 = _T_73 | out_live_in_fire_R_8_0; // @[LoopBlock.scala 722:57]
  assign _T_74 = io_OutLiveIn_field9_0_ready & io_OutLiveIn_field9_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_96 = _T_74 ? 1'h0 : out_live_in_valid_R_9_0; // @[LoopBlock.scala 722:57]
  assign _GEN_97 = _T_74 | out_live_in_fire_R_9_0; // @[LoopBlock.scala 722:57]
  assign _T_75 = io_OutLiveIn_field10_0_ready & io_OutLiveIn_field10_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_98 = _T_75 ? 1'h0 : out_live_in_valid_R_10_0; // @[LoopBlock.scala 722:57]
  assign _GEN_99 = _T_75 | out_live_in_fire_R_10_0; // @[LoopBlock.scala 722:57]
  assign _T_76 = io_OutLiveIn_field11_0_ready & io_OutLiveIn_field11_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_100 = _T_76 ? 1'h0 : out_live_in_valid_R_11_0; // @[LoopBlock.scala 722:57]
  assign _GEN_101 = _T_76 | out_live_in_fire_R_11_0; // @[LoopBlock.scala 722:57]
  assign _T_77 = io_OutLiveIn_field12_0_ready & io_OutLiveIn_field12_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_102 = _T_77 ? 1'h0 : out_live_in_valid_R_12_0; // @[LoopBlock.scala 722:57]
  assign _GEN_103 = _T_77 | out_live_in_fire_R_12_0; // @[LoopBlock.scala 722:57]
  assign _T_78 = io_CarryDepenOut_field0_0_ready & io_CarryDepenOut_field0_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_104 = _T_78 ? 1'h0 : out_carry_out_valid_R_0_0; // @[LoopBlock.scala 742:61]
  assign _T_79 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_80 = in_live_in_valid_R_0 & in_live_in_valid_R_1; // @[LoopBlock.scala 765:35]
  assign _T_81 = _T_80 & in_live_in_valid_R_2; // @[LoopBlock.scala 765:35]
  assign _T_82 = _T_81 & in_live_in_valid_R_3; // @[LoopBlock.scala 765:35]
  assign _T_83 = _T_82 & in_live_in_valid_R_4; // @[LoopBlock.scala 765:35]
  assign _T_84 = _T_83 & in_live_in_valid_R_5; // @[LoopBlock.scala 765:35]
  assign _T_85 = _T_84 & in_live_in_valid_R_6; // @[LoopBlock.scala 765:35]
  assign _T_86 = _T_85 & in_live_in_valid_R_7; // @[LoopBlock.scala 765:35]
  assign _T_87 = _T_86 & in_live_in_valid_R_8; // @[LoopBlock.scala 765:35]
  assign _T_88 = _T_87 & in_live_in_valid_R_9; // @[LoopBlock.scala 765:35]
  assign _T_89 = _T_88 & in_live_in_valid_R_10; // @[LoopBlock.scala 765:35]
  assign _T_90 = _T_89 & in_live_in_valid_R_11; // @[LoopBlock.scala 765:35]
  assign _T_91 = _T_90 & in_live_in_valid_R_12; // @[LoopBlock.scala 765:35]
  assign _T_92 = _T_91 & enable_valid_R; // @[LoopBlock.scala 869:28]
  assign _GEN_106 = enable_R_control | _GEN_70; // @[LoopBlock.scala 870:26]
  assign _GEN_107 = enable_R_control | _GEN_72; // @[LoopBlock.scala 870:26]
  assign _GEN_108 = enable_R_control | _GEN_74; // @[LoopBlock.scala 870:26]
  assign _GEN_109 = enable_R_control | _GEN_76; // @[LoopBlock.scala 870:26]
  assign _GEN_110 = enable_R_control | _GEN_78; // @[LoopBlock.scala 870:26]
  assign _GEN_111 = enable_R_control | _GEN_80; // @[LoopBlock.scala 870:26]
  assign _GEN_112 = enable_R_control | _GEN_82; // @[LoopBlock.scala 870:26]
  assign _GEN_113 = enable_R_control | _GEN_84; // @[LoopBlock.scala 870:26]
  assign _GEN_114 = enable_R_control | _GEN_86; // @[LoopBlock.scala 870:26]
  assign _GEN_115 = enable_R_control | _GEN_88; // @[LoopBlock.scala 870:26]
  assign _GEN_116 = enable_R_control | _GEN_90; // @[LoopBlock.scala 870:26]
  assign _GEN_117 = enable_R_control | _GEN_92; // @[LoopBlock.scala 870:26]
  assign _GEN_118 = enable_R_control | _GEN_94; // @[LoopBlock.scala 870:26]
  assign _GEN_119 = enable_R_control | _GEN_96; // @[LoopBlock.scala 870:26]
  assign _GEN_120 = enable_R_control | _GEN_98; // @[LoopBlock.scala 870:26]
  assign _GEN_121 = enable_R_control | _GEN_100; // @[LoopBlock.scala 870:26]
  assign _GEN_122 = enable_R_control | _GEN_102; // @[LoopBlock.scala 870:26]
  assign _GEN_123 = enable_R_control | _GEN_104; // @[LoopBlock.scala 870:26]
  assign _GEN_124 = enable_R_control | active_loop_start_R_control; // @[LoopBlock.scala 870:26]
  assign _GEN_126 = enable_R_control | _GEN_66; // @[LoopBlock.scala 870:26]
  assign _GEN_129 = enable_R_control | _GEN_67; // @[LoopBlock.scala 870:26]
  assign _GEN_131 = enable_R_control & loop_exit_R_0_control; // @[LoopBlock.scala 870:26]
  assign _T_96 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_97 = loop_back_valid_R_0 & loop_finish_valid_R_0; // @[LoopBlock.scala 898:30]
  assign _T_99 = out_live_in_fire_R_0_0 & out_live_in_fire_R_0_1; // @[LoopBlock.scala 825:65]
  assign _T_100 = _T_99 & out_live_in_fire_R_0_2; // @[LoopBlock.scala 825:65]
  assign _T_101 = out_live_in_fire_R_1_0 & out_live_in_fire_R_1_1; // @[LoopBlock.scala 825:65]
  assign _T_102 = _T_101 & out_live_in_fire_R_1_2; // @[LoopBlock.scala 825:65]
  assign _T_103 = _T_100 & _T_102; // @[LoopBlock.scala 828:26]
  assign _T_104 = _T_103 & out_live_in_fire_R_2_0; // @[LoopBlock.scala 828:26]
  assign _T_105 = _T_104 & out_live_in_fire_R_3_0; // @[LoopBlock.scala 828:26]
  assign _T_106 = _T_105 & out_live_in_fire_R_4_0; // @[LoopBlock.scala 828:26]
  assign _T_107 = _T_106 & out_live_in_fire_R_5_0; // @[LoopBlock.scala 828:26]
  assign _T_108 = _T_107 & out_live_in_fire_R_6_0; // @[LoopBlock.scala 828:26]
  assign _T_109 = _T_108 & out_live_in_fire_R_7_0; // @[LoopBlock.scala 828:26]
  assign _T_110 = _T_109 & out_live_in_fire_R_8_0; // @[LoopBlock.scala 828:26]
  assign _T_111 = _T_110 & out_live_in_fire_R_9_0; // @[LoopBlock.scala 828:26]
  assign _T_112 = _T_111 & out_live_in_fire_R_10_0; // @[LoopBlock.scala 828:26]
  assign _T_113 = _T_112 & out_live_in_fire_R_11_0; // @[LoopBlock.scala 828:26]
  assign _T_114 = _T_113 & out_live_in_fire_R_12_0; // @[LoopBlock.scala 828:26]
  assign _T_115 = _T_97 & _T_114; // @[LoopBlock.scala 899:29]
  assign _T_122 = $unsigned(reset); // @[LoopBlock.scala 932:19]
  assign _T_123 = _T_122 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_162 = loop_finish_R_0_control | _GEN_68; // @[LoopBlock.scala 936:64]
  assign _GEN_165 = loop_finish_R_0_control ? 1'h0 : active_loop_back_R_control; // @[LoopBlock.scala 936:64]
  assign _GEN_167 = loop_finish_R_0_control | loop_exit_R_0_control; // @[LoopBlock.scala 936:64]
  assign _GEN_172 = loop_back_R_0_control | _GEN_66; // @[LoopBlock.scala 903:56]
  assign _GEN_173 = loop_back_R_0_control | _GEN_165; // @[LoopBlock.scala 903:56]
  assign _GEN_175 = loop_back_R_0_control | _GEN_67; // @[LoopBlock.scala 903:56]
  assign _GEN_194 = loop_back_R_0_control | _GEN_70; // @[LoopBlock.scala 903:56]
  assign _GEN_195 = loop_back_R_0_control | _GEN_72; // @[LoopBlock.scala 903:56]
  assign _GEN_196 = loop_back_R_0_control | _GEN_74; // @[LoopBlock.scala 903:56]
  assign _GEN_197 = loop_back_R_0_control | _GEN_76; // @[LoopBlock.scala 903:56]
  assign _GEN_198 = loop_back_R_0_control | _GEN_78; // @[LoopBlock.scala 903:56]
  assign _GEN_199 = loop_back_R_0_control | _GEN_80; // @[LoopBlock.scala 903:56]
  assign _GEN_200 = loop_back_R_0_control | _GEN_82; // @[LoopBlock.scala 903:56]
  assign _GEN_201 = loop_back_R_0_control | _GEN_84; // @[LoopBlock.scala 903:56]
  assign _GEN_202 = loop_back_R_0_control | _GEN_86; // @[LoopBlock.scala 903:56]
  assign _GEN_203 = loop_back_R_0_control | _GEN_88; // @[LoopBlock.scala 903:56]
  assign _GEN_204 = loop_back_R_0_control | _GEN_90; // @[LoopBlock.scala 903:56]
  assign _GEN_205 = loop_back_R_0_control | _GEN_92; // @[LoopBlock.scala 903:56]
  assign _GEN_206 = loop_back_R_0_control | _GEN_94; // @[LoopBlock.scala 903:56]
  assign _GEN_207 = loop_back_R_0_control | _GEN_96; // @[LoopBlock.scala 903:56]
  assign _GEN_208 = loop_back_R_0_control | _GEN_98; // @[LoopBlock.scala 903:56]
  assign _GEN_209 = loop_back_R_0_control | _GEN_100; // @[LoopBlock.scala 903:56]
  assign _GEN_210 = loop_back_R_0_control | _GEN_102; // @[LoopBlock.scala 903:56]
  assign _GEN_211 = loop_back_R_0_control | _GEN_104; // @[LoopBlock.scala 903:56]
  assign _T_131 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[LoopBlock.scala 595:19]
  assign io_InLiveIn_0_ready = ~ in_live_in_valid_R_0; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_1_ready = ~ in_live_in_valid_R_1; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_2_ready = ~ in_live_in_valid_R_2; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_3_ready = ~ in_live_in_valid_R_3; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_4_ready = ~ in_live_in_valid_R_4; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_5_ready = ~ in_live_in_valid_R_5; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_6_ready = ~ in_live_in_valid_R_6; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_7_ready = ~ in_live_in_valid_R_7; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_8_ready = ~ in_live_in_valid_R_8; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_9_ready = ~ in_live_in_valid_R_9; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_10_ready = ~ in_live_in_valid_R_10; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_11_ready = ~ in_live_in_valid_R_11; // @[LoopBlock.scala 622:26]
  assign io_InLiveIn_12_ready = ~ in_live_in_valid_R_12; // @[LoopBlock.scala 622:26]
  assign io_OutLiveIn_field12_0_valid = out_live_in_valid_R_12_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field12_0_bits_predicate = in_live_in_R_12_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field12_0_bits_taskID = in_live_in_R_12_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field12_0_bits_data = in_live_in_R_12_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field11_0_valid = out_live_in_valid_R_11_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field11_0_bits_predicate = in_live_in_R_11_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field11_0_bits_taskID = in_live_in_R_11_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field11_0_bits_data = in_live_in_R_11_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_0_valid = out_live_in_valid_R_10_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field10_0_bits_predicate = in_live_in_R_10_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_0_bits_taskID = in_live_in_R_10_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field10_0_bits_data = in_live_in_R_10_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field9_0_valid = out_live_in_valid_R_9_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field9_0_bits_predicate = in_live_in_R_9_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field9_0_bits_taskID = in_live_in_R_9_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field9_0_bits_data = in_live_in_R_9_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_valid = out_live_in_valid_R_8_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field8_0_bits_predicate = in_live_in_R_8_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_bits_taskID = in_live_in_R_8_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field8_0_bits_data = in_live_in_R_8_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_valid = out_live_in_valid_R_7_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field7_0_bits_predicate = in_live_in_R_7_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_bits_taskID = in_live_in_R_7_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field7_0_bits_data = in_live_in_R_7_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_valid = out_live_in_valid_R_6_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field6_0_bits_predicate = in_live_in_R_6_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_bits_taskID = in_live_in_R_6_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field6_0_bits_data = in_live_in_R_6_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_0_valid = out_live_in_valid_R_5_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field5_0_bits_predicate = in_live_in_R_5_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_0_bits_taskID = in_live_in_R_5_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field5_0_bits_data = in_live_in_R_5_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_valid = out_live_in_valid_R_4_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field4_0_bits_taskID = in_live_in_R_4_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field4_0_bits_data = in_live_in_R_4_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_valid = out_live_in_valid_R_3_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field3_0_bits_predicate = in_live_in_R_3_predicate; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_bits_taskID = in_live_in_R_3_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field3_0_bits_data = in_live_in_R_3_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_valid = out_live_in_valid_R_2_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field2_0_bits_taskID = in_live_in_R_2_taskID; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field2_0_bits_data = in_live_in_R_2_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_0_valid = out_live_in_valid_R_1_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_0_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_1_valid = out_live_in_valid_R_1_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_1_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field1_2_valid = out_live_in_valid_R_1_2; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field1_2_bits_data = in_live_in_R_1_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_0_valid = out_live_in_valid_R_0_0; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_0_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_1_valid = out_live_in_valid_R_0_1; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_1_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_OutLiveIn_field0_2_valid = out_live_in_valid_R_0_2; // @[LoopBlock.scala 665:50]
  assign io_OutLiveIn_field0_2_bits_data = in_live_in_R_0_data; // @[LoopBlock.scala 664:49]
  assign io_activate_loop_start_valid = active_loop_start_valid_R; // @[LoopBlock.scala 689:32]
  assign io_activate_loop_start_bits_taskID = active_loop_start_R_taskID; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_start_bits_control = active_loop_start_R_control; // @[LoopBlock.scala 688:31]
  assign io_activate_loop_back_valid = active_loop_back_valid_R; // @[LoopBlock.scala 692:31]
  assign io_activate_loop_back_bits_taskID = active_loop_back_R_taskID; // @[LoopBlock.scala 691:30]
  assign io_activate_loop_back_bits_control = active_loop_back_R_control; // @[LoopBlock.scala 691:30]
  assign io_loopBack_0_ready = ~ loop_back_valid_R_0; // @[LoopBlock.scala 602:26]
  assign io_loopFinish_0_ready = ~ loop_finish_valid_R_0; // @[LoopBlock.scala 611:28]
  assign io_CarryDepenIn_0_ready = ~ in_carry_in_valid_R_0; // @[LoopBlock.scala 640:30]
  assign io_CarryDepenOut_field0_0_valid = out_carry_out_valid_R_0_0; // @[LoopBlock.scala 681:54]
  assign io_CarryDepenOut_field0_0_bits_taskID = in_carry_in_R_0_taskID; // @[LoopBlock.scala 680:53]
  assign io_CarryDepenOut_field0_0_bits_data = in_carry_in_R_0_data; // @[LoopBlock.scala 680:53]
  assign io_loopExit_0_valid = loop_exit_valid_R_0; // @[LoopBlock.scala 696:26]
  assign io_loopExit_0_bits_taskID = loop_exit_R_0_taskID; // @[LoopBlock.scala 695:25]
  assign io_loopExit_0_bits_control = loop_exit_R_0_control; // @[LoopBlock.scala 695:25]
  assign _GEN_618 = _T_79 == 1'h0; // @[LoopBlock.scala 932:19]
  assign _GEN_619 = _GEN_618 & _T_96; // @[LoopBlock.scala 932:19]
  assign _GEN_620 = _GEN_619 & _T_115; // @[LoopBlock.scala 932:19]
  assign _GEN_621 = _GEN_620 & loop_back_R_0_control; // @[LoopBlock.scala 932:19]
  assign _GEN_625 = loop_back_R_0_control == 1'h0; // @[LoopBlock.scala 950:19]
  assign _GEN_626 = _GEN_620 & _GEN_625; // @[LoopBlock.scala 950:19]
  assign _GEN_627 = _GEN_626 & loop_finish_R_0_control; // @[LoopBlock.scala 950:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_valid_R = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  loop_back_R_0_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  loop_back_R_0_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  loop_back_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  loop_finish_R_0_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  loop_finish_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  in_live_in_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  in_live_in_R_1_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  in_live_in_R_2_taskID = _RAND_11[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  in_live_in_R_2_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  in_live_in_R_3_predicate = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  in_live_in_R_3_taskID = _RAND_14[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  in_live_in_R_3_data = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  in_live_in_R_4_taskID = _RAND_16[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  in_live_in_R_4_data = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  in_live_in_R_5_predicate = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  in_live_in_R_5_taskID = _RAND_19[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  in_live_in_R_5_data = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  in_live_in_R_6_predicate = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  in_live_in_R_6_taskID = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  in_live_in_R_6_data = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  in_live_in_R_7_predicate = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  in_live_in_R_7_taskID = _RAND_25[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  in_live_in_R_7_data = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  in_live_in_R_8_predicate = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  in_live_in_R_8_taskID = _RAND_28[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  in_live_in_R_8_data = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  in_live_in_R_9_predicate = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  in_live_in_R_9_taskID = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  in_live_in_R_9_data = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  in_live_in_R_10_predicate = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  in_live_in_R_10_taskID = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  in_live_in_R_10_data = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  in_live_in_R_11_predicate = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  in_live_in_R_11_taskID = _RAND_37[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  in_live_in_R_11_data = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  in_live_in_R_12_predicate = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  in_live_in_R_12_taskID = _RAND_40[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  in_live_in_R_12_data = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  in_live_in_valid_R_0 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  in_live_in_valid_R_1 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  in_live_in_valid_R_2 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  in_live_in_valid_R_3 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  in_live_in_valid_R_4 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  in_live_in_valid_R_5 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  in_live_in_valid_R_6 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  in_live_in_valid_R_7 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  in_live_in_valid_R_8 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  in_live_in_valid_R_9 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  in_live_in_valid_R_10 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  in_live_in_valid_R_11 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  in_live_in_valid_R_12 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  in_carry_in_R_0_taskID = _RAND_55[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  in_carry_in_R_0_data = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  in_carry_in_valid_R_0 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  out_live_in_valid_R_0_0 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  out_live_in_valid_R_0_1 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  out_live_in_valid_R_0_2 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  out_live_in_valid_R_1_0 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  out_live_in_valid_R_1_1 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  out_live_in_valid_R_1_2 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  out_live_in_valid_R_2_0 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  out_live_in_valid_R_3_0 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  out_live_in_valid_R_4_0 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  out_live_in_valid_R_5_0 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  out_live_in_valid_R_6_0 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  out_live_in_valid_R_7_0 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  out_live_in_valid_R_8_0 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  out_live_in_valid_R_9_0 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  out_live_in_valid_R_10_0 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  out_live_in_valid_R_11_0 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  out_live_in_valid_R_12_0 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  out_live_in_fire_R_0_0 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  out_live_in_fire_R_0_1 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  out_live_in_fire_R_0_2 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  out_live_in_fire_R_1_0 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  out_live_in_fire_R_1_1 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  out_live_in_fire_R_1_2 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  out_live_in_fire_R_2_0 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  out_live_in_fire_R_3_0 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  out_live_in_fire_R_4_0 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  out_live_in_fire_R_5_0 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  out_live_in_fire_R_6_0 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  out_live_in_fire_R_7_0 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  out_live_in_fire_R_8_0 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  out_live_in_fire_R_9_0 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  out_live_in_fire_R_10_0 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  out_live_in_fire_R_11_0 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  out_live_in_fire_R_12_0 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  out_carry_out_valid_R_0_0 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  active_loop_start_R_taskID = _RAND_93[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  active_loop_start_R_control = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  active_loop_start_valid_R = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  active_loop_back_R_taskID = _RAND_96[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  active_loop_back_R_control = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  active_loop_back_valid_R = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  loop_exit_R_0_taskID = _RAND_99[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  loop_exit_R_0_control = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  loop_exit_valid_R_0 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  loop_exit_fire_R_0 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  state = _RAND_103[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_25) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_25) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              enable_R_taskID <= 5'h0;
            end else begin
              if (_T_25) begin
                enable_R_taskID <= io_enable_bits_taskID;
              end
            end
          end else begin
            if (_T_25) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_25) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_96) begin
          if (_T_25) begin
            enable_R_control <= io_enable_bits_control;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_25) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_25) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_79) begin
        enable_valid_R <= _GEN_3;
      end else begin
        if (_T_96) begin
          enable_valid_R <= _GEN_3;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_3;
            end
          end else begin
            enable_valid_R <= _GEN_3;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_27) begin
          loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_27) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            if (_T_27) begin
              loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
            end
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_taskID <= 5'h0;
            end else begin
              if (_T_27) begin
                loop_back_R_0_taskID <= io_loopBack_0_bits_taskID;
              end
            end
          end else begin
            loop_back_R_0_taskID <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      loop_back_R_0_control <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_27) begin
          loop_back_R_0_control <= io_loopBack_0_bits_control;
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_27) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            if (_T_27) begin
              loop_back_R_0_control <= io_loopBack_0_bits_control;
            end
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              loop_back_R_0_control <= 1'h0;
            end else begin
              if (_T_27) begin
                loop_back_R_0_control <= io_loopBack_0_bits_control;
              end
            end
          end else begin
            loop_back_R_0_control <= _GEN_4;
          end
        end
      end
    end
    if (reset) begin
      loop_back_valid_R_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        loop_back_valid_R_0 <= _GEN_6;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              loop_back_valid_R_0 <= 1'h0;
            end else begin
              loop_back_valid_R_0 <= _GEN_6;
            end
          end else begin
            loop_back_valid_R_0 <= _GEN_6;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_R_0_control <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_29) begin
          loop_finish_R_0_control <= io_loopFinish_0_bits_control;
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_29) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            if (_T_29) begin
              loop_finish_R_0_control <= io_loopFinish_0_bits_control;
            end
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_R_0_control <= 1'h0;
            end else begin
              if (_T_29) begin
                loop_finish_R_0_control <= io_loopFinish_0_bits_control;
              end
            end
          end else begin
            loop_finish_R_0_control <= _GEN_7;
          end
        end
      end
    end
    if (reset) begin
      loop_finish_valid_R_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        loop_finish_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              loop_finish_valid_R_0 <= 1'h0;
            end else begin
              loop_finish_valid_R_0 <= _GEN_9;
            end
          end else begin
            loop_finish_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_0_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_31) begin
          in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_31) begin
            in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_0_data <= 32'h0;
            end else begin
              if (_T_31) begin
                in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
              end
            end
          end else begin
            if (_T_31) begin
              in_live_in_R_0_data <= io_InLiveIn_0_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_1_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_33) begin
          in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_33) begin
            in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_1_data <= 32'h0;
            end else begin
              if (_T_33) begin
                in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
              end
            end
          end else begin
            if (_T_33) begin
              in_live_in_R_1_data <= io_InLiveIn_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_35) begin
          in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_35) begin
            in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_taskID <= 5'h0;
            end else begin
              if (_T_35) begin
                in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
              end
            end
          end else begin
            if (_T_35) begin
              in_live_in_R_2_taskID <= io_InLiveIn_2_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_2_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_35) begin
          in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_35) begin
            in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_2_data <= 32'h0;
            end else begin
              if (_T_35) begin
                in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
              end
            end
          end else begin
            if (_T_35) begin
              in_live_in_R_2_data <= io_InLiveIn_2_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_predicate <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_37) begin
          in_live_in_R_3_predicate <= io_InLiveIn_3_bits_predicate;
        end
      end else begin
        if (_T_96) begin
          if (_T_37) begin
            in_live_in_R_3_predicate <= io_InLiveIn_3_bits_predicate;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_predicate <= 1'h0;
            end else begin
              if (_T_37) begin
                in_live_in_R_3_predicate <= io_InLiveIn_3_bits_predicate;
              end
            end
          end else begin
            if (_T_37) begin
              in_live_in_R_3_predicate <= io_InLiveIn_3_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_37) begin
          in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_37) begin
            in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_taskID <= 5'h0;
            end else begin
              if (_T_37) begin
                in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
              end
            end
          end else begin
            if (_T_37) begin
              in_live_in_R_3_taskID <= io_InLiveIn_3_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_3_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_37) begin
          in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_37) begin
            in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_3_data <= 32'h0;
            end else begin
              if (_T_37) begin
                in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
              end
            end
          end else begin
            if (_T_37) begin
              in_live_in_R_3_data <= io_InLiveIn_3_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_39) begin
          in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_39) begin
            in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_taskID <= 5'h0;
            end else begin
              if (_T_39) begin
                in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
              end
            end
          end else begin
            if (_T_39) begin
              in_live_in_R_4_taskID <= io_InLiveIn_4_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_4_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_39) begin
          in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_39) begin
            in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_4_data <= 32'h0;
            end else begin
              if (_T_39) begin
                in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
              end
            end
          end else begin
            if (_T_39) begin
              in_live_in_R_4_data <= io_InLiveIn_4_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_predicate <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_41) begin
          in_live_in_R_5_predicate <= io_InLiveIn_5_bits_predicate;
        end
      end else begin
        if (_T_96) begin
          if (_T_41) begin
            in_live_in_R_5_predicate <= io_InLiveIn_5_bits_predicate;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_predicate <= 1'h0;
            end else begin
              if (_T_41) begin
                in_live_in_R_5_predicate <= io_InLiveIn_5_bits_predicate;
              end
            end
          end else begin
            if (_T_41) begin
              in_live_in_R_5_predicate <= io_InLiveIn_5_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_41) begin
          in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_41) begin
            in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_taskID <= 5'h0;
            end else begin
              if (_T_41) begin
                in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
              end
            end
          end else begin
            if (_T_41) begin
              in_live_in_R_5_taskID <= io_InLiveIn_5_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_5_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_41) begin
          in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_41) begin
            in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_5_data <= 32'h0;
            end else begin
              if (_T_41) begin
                in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
              end
            end
          end else begin
            if (_T_41) begin
              in_live_in_R_5_data <= io_InLiveIn_5_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_predicate <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_43) begin
          in_live_in_R_6_predicate <= io_InLiveIn_6_bits_predicate;
        end
      end else begin
        if (_T_96) begin
          if (_T_43) begin
            in_live_in_R_6_predicate <= io_InLiveIn_6_bits_predicate;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_predicate <= 1'h0;
            end else begin
              if (_T_43) begin
                in_live_in_R_6_predicate <= io_InLiveIn_6_bits_predicate;
              end
            end
          end else begin
            if (_T_43) begin
              in_live_in_R_6_predicate <= io_InLiveIn_6_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_43) begin
          in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_43) begin
            in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_taskID <= 5'h0;
            end else begin
              if (_T_43) begin
                in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
              end
            end
          end else begin
            if (_T_43) begin
              in_live_in_R_6_taskID <= io_InLiveIn_6_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_6_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_43) begin
          in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_43) begin
            in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_6_data <= 32'h0;
            end else begin
              if (_T_43) begin
                in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
              end
            end
          end else begin
            if (_T_43) begin
              in_live_in_R_6_data <= io_InLiveIn_6_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_predicate <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_45) begin
          in_live_in_R_7_predicate <= io_InLiveIn_7_bits_predicate;
        end
      end else begin
        if (_T_96) begin
          if (_T_45) begin
            in_live_in_R_7_predicate <= io_InLiveIn_7_bits_predicate;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_predicate <= 1'h0;
            end else begin
              if (_T_45) begin
                in_live_in_R_7_predicate <= io_InLiveIn_7_bits_predicate;
              end
            end
          end else begin
            if (_T_45) begin
              in_live_in_R_7_predicate <= io_InLiveIn_7_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_45) begin
          in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_45) begin
            in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_taskID <= 5'h0;
            end else begin
              if (_T_45) begin
                in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
              end
            end
          end else begin
            if (_T_45) begin
              in_live_in_R_7_taskID <= io_InLiveIn_7_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_7_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_45) begin
          in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_45) begin
            in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_7_data <= 32'h0;
            end else begin
              if (_T_45) begin
                in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
              end
            end
          end else begin
            if (_T_45) begin
              in_live_in_R_7_data <= io_InLiveIn_7_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_predicate <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_47) begin
          in_live_in_R_8_predicate <= io_InLiveIn_8_bits_predicate;
        end
      end else begin
        if (_T_96) begin
          if (_T_47) begin
            in_live_in_R_8_predicate <= io_InLiveIn_8_bits_predicate;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_predicate <= 1'h0;
            end else begin
              if (_T_47) begin
                in_live_in_R_8_predicate <= io_InLiveIn_8_bits_predicate;
              end
            end
          end else begin
            if (_T_47) begin
              in_live_in_R_8_predicate <= io_InLiveIn_8_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_47) begin
          in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_47) begin
            in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_taskID <= 5'h0;
            end else begin
              if (_T_47) begin
                in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
              end
            end
          end else begin
            if (_T_47) begin
              in_live_in_R_8_taskID <= io_InLiveIn_8_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_8_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_47) begin
          in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_47) begin
            in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_8_data <= 32'h0;
            end else begin
              if (_T_47) begin
                in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
              end
            end
          end else begin
            if (_T_47) begin
              in_live_in_R_8_data <= io_InLiveIn_8_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_9_predicate <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_49) begin
          in_live_in_R_9_predicate <= io_InLiveIn_9_bits_predicate;
        end
      end else begin
        if (_T_96) begin
          if (_T_49) begin
            in_live_in_R_9_predicate <= io_InLiveIn_9_bits_predicate;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_9_predicate <= 1'h0;
            end else begin
              if (_T_49) begin
                in_live_in_R_9_predicate <= io_InLiveIn_9_bits_predicate;
              end
            end
          end else begin
            if (_T_49) begin
              in_live_in_R_9_predicate <= io_InLiveIn_9_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_9_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_49) begin
          in_live_in_R_9_taskID <= io_InLiveIn_9_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_49) begin
            in_live_in_R_9_taskID <= io_InLiveIn_9_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_9_taskID <= 5'h0;
            end else begin
              if (_T_49) begin
                in_live_in_R_9_taskID <= io_InLiveIn_9_bits_taskID;
              end
            end
          end else begin
            if (_T_49) begin
              in_live_in_R_9_taskID <= io_InLiveIn_9_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_9_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_49) begin
          in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_49) begin
            in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_9_data <= 32'h0;
            end else begin
              if (_T_49) begin
                in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
              end
            end
          end else begin
            if (_T_49) begin
              in_live_in_R_9_data <= io_InLiveIn_9_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_10_predicate <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_51) begin
          in_live_in_R_10_predicate <= io_InLiveIn_10_bits_predicate;
        end
      end else begin
        if (_T_96) begin
          if (_T_51) begin
            in_live_in_R_10_predicate <= io_InLiveIn_10_bits_predicate;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_10_predicate <= 1'h0;
            end else begin
              if (_T_51) begin
                in_live_in_R_10_predicate <= io_InLiveIn_10_bits_predicate;
              end
            end
          end else begin
            if (_T_51) begin
              in_live_in_R_10_predicate <= io_InLiveIn_10_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_10_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_51) begin
          in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_51) begin
            in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_10_taskID <= 5'h0;
            end else begin
              if (_T_51) begin
                in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
              end
            end
          end else begin
            if (_T_51) begin
              in_live_in_R_10_taskID <= io_InLiveIn_10_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_10_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_51) begin
          in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_51) begin
            in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_10_data <= 32'h0;
            end else begin
              if (_T_51) begin
                in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
              end
            end
          end else begin
            if (_T_51) begin
              in_live_in_R_10_data <= io_InLiveIn_10_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_11_predicate <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_53) begin
          in_live_in_R_11_predicate <= io_InLiveIn_11_bits_predicate;
        end
      end else begin
        if (_T_96) begin
          if (_T_53) begin
            in_live_in_R_11_predicate <= io_InLiveIn_11_bits_predicate;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_11_predicate <= 1'h0;
            end else begin
              if (_T_53) begin
                in_live_in_R_11_predicate <= io_InLiveIn_11_bits_predicate;
              end
            end
          end else begin
            if (_T_53) begin
              in_live_in_R_11_predicate <= io_InLiveIn_11_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_11_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_53) begin
          in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_53) begin
            in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_11_taskID <= 5'h0;
            end else begin
              if (_T_53) begin
                in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
              end
            end
          end else begin
            if (_T_53) begin
              in_live_in_R_11_taskID <= io_InLiveIn_11_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_11_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_53) begin
          in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_53) begin
            in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_11_data <= 32'h0;
            end else begin
              if (_T_53) begin
                in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
              end
            end
          end else begin
            if (_T_53) begin
              in_live_in_R_11_data <= io_InLiveIn_11_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_12_predicate <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_55) begin
          in_live_in_R_12_predicate <= io_InLiveIn_12_bits_predicate;
        end
      end else begin
        if (_T_96) begin
          if (_T_55) begin
            in_live_in_R_12_predicate <= io_InLiveIn_12_bits_predicate;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_12_predicate <= 1'h0;
            end else begin
              if (_T_55) begin
                in_live_in_R_12_predicate <= io_InLiveIn_12_bits_predicate;
              end
            end
          end else begin
            if (_T_55) begin
              in_live_in_R_12_predicate <= io_InLiveIn_12_bits_predicate;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_12_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_55) begin
          in_live_in_R_12_taskID <= io_InLiveIn_12_bits_taskID;
        end
      end else begin
        if (_T_96) begin
          if (_T_55) begin
            in_live_in_R_12_taskID <= io_InLiveIn_12_bits_taskID;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_12_taskID <= 5'h0;
            end else begin
              if (_T_55) begin
                in_live_in_R_12_taskID <= io_InLiveIn_12_bits_taskID;
              end
            end
          end else begin
            if (_T_55) begin
              in_live_in_R_12_taskID <= io_InLiveIn_12_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_R_12_data <= 32'h0;
    end else begin
      if (_T_79) begin
        if (_T_55) begin
          in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
        end
      end else begin
        if (_T_96) begin
          if (_T_55) begin
            in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_R_12_data <= 32'h0;
            end else begin
              if (_T_55) begin
                in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
              end
            end
          end else begin
            if (_T_55) begin
              in_live_in_R_12_data <= io_InLiveIn_12_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_0 <= _GEN_13;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_0 <= _GEN_13;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_0 <= 1'h0;
            end else begin
              in_live_in_valid_R_0 <= _GEN_13;
            end
          end else begin
            in_live_in_valid_R_0 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_1 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_1 <= _GEN_17;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_1 <= _GEN_17;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_1 <= 1'h0;
            end else begin
              in_live_in_valid_R_1 <= _GEN_17;
            end
          end else begin
            in_live_in_valid_R_1 <= _GEN_17;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_2 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_2 <= _GEN_21;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_2 <= _GEN_21;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_2 <= 1'h0;
            end else begin
              in_live_in_valid_R_2 <= _GEN_21;
            end
          end else begin
            in_live_in_valid_R_2 <= _GEN_21;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_3 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_3 <= _GEN_25;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_3 <= _GEN_25;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_3 <= 1'h0;
            end else begin
              in_live_in_valid_R_3 <= _GEN_25;
            end
          end else begin
            in_live_in_valid_R_3 <= _GEN_25;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_4 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_4 <= _GEN_29;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_4 <= _GEN_29;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_4 <= 1'h0;
            end else begin
              in_live_in_valid_R_4 <= _GEN_29;
            end
          end else begin
            in_live_in_valid_R_4 <= _GEN_29;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_5 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_5 <= _GEN_33;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_5 <= _GEN_33;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_5 <= 1'h0;
            end else begin
              in_live_in_valid_R_5 <= _GEN_33;
            end
          end else begin
            in_live_in_valid_R_5 <= _GEN_33;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_6 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_6 <= _GEN_37;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_6 <= _GEN_37;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_6 <= 1'h0;
            end else begin
              in_live_in_valid_R_6 <= _GEN_37;
            end
          end else begin
            in_live_in_valid_R_6 <= _GEN_37;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_7 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_7 <= _GEN_41;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_7 <= _GEN_41;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_7 <= 1'h0;
            end else begin
              in_live_in_valid_R_7 <= _GEN_41;
            end
          end else begin
            in_live_in_valid_R_7 <= _GEN_41;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_8 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_8 <= _GEN_45;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_8 <= _GEN_45;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_8 <= 1'h0;
            end else begin
              in_live_in_valid_R_8 <= _GEN_45;
            end
          end else begin
            in_live_in_valid_R_8 <= _GEN_45;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_9 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_9 <= _GEN_49;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_9 <= _GEN_49;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_9 <= 1'h0;
            end else begin
              in_live_in_valid_R_9 <= _GEN_49;
            end
          end else begin
            in_live_in_valid_R_9 <= _GEN_49;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_10 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_10 <= _GEN_53;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_10 <= _GEN_53;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_10 <= 1'h0;
            end else begin
              in_live_in_valid_R_10 <= _GEN_53;
            end
          end else begin
            in_live_in_valid_R_10 <= _GEN_53;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_11 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_11 <= _GEN_57;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_11 <= _GEN_57;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_11 <= 1'h0;
            end else begin
              in_live_in_valid_R_11 <= _GEN_57;
            end
          end else begin
            in_live_in_valid_R_11 <= _GEN_57;
          end
        end
      end
    end
    if (reset) begin
      in_live_in_valid_R_12 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_live_in_valid_R_12 <= _GEN_61;
      end else begin
        if (_T_96) begin
          in_live_in_valid_R_12 <= _GEN_61;
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_live_in_valid_R_12 <= 1'h0;
            end else begin
              in_live_in_valid_R_12 <= _GEN_61;
            end
          end else begin
            in_live_in_valid_R_12 <= _GEN_61;
          end
        end
      end
    end
    if (reset) begin
      in_carry_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_57) begin
        in_carry_in_R_0_taskID <= io_CarryDepenIn_0_bits_taskID;
      end
    end
    if (reset) begin
      in_carry_in_R_0_data <= 32'h0;
    end else begin
      if (_T_57) begin
        in_carry_in_R_0_data <= io_CarryDepenIn_0_bits_data;
      end
    end
    if (reset) begin
      in_carry_in_valid_R_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        in_carry_in_valid_R_0 <= _GEN_65;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_65;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_65;
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              in_carry_in_valid_R_0 <= 1'h0;
            end else begin
              in_carry_in_valid_R_0 <= _GEN_65;
            end
          end else begin
            in_carry_in_valid_R_0 <= _GEN_65;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_0_0 <= _GEN_106;
        end else begin
          if (_T_61) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_0_0 <= _GEN_194;
          end else begin
            if (_T_61) begin
              out_live_in_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_61) begin
            out_live_in_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_1 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_0_1 <= _GEN_107;
        end else begin
          if (_T_62) begin
            out_live_in_valid_R_0_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_0_1 <= _GEN_195;
          end else begin
            if (_T_62) begin
              out_live_in_valid_R_0_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_62) begin
            out_live_in_valid_R_0_1 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_0_2 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_0_2 <= _GEN_108;
        end else begin
          if (_T_63) begin
            out_live_in_valid_R_0_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_0_2 <= _GEN_196;
          end else begin
            if (_T_63) begin
              out_live_in_valid_R_0_2 <= 1'h0;
            end
          end
        end else begin
          if (_T_63) begin
            out_live_in_valid_R_0_2 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_1_0 <= _GEN_109;
        end else begin
          if (_T_64) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_1_0 <= _GEN_197;
          end else begin
            if (_T_64) begin
              out_live_in_valid_R_1_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_64) begin
            out_live_in_valid_R_1_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_1 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_1_1 <= _GEN_110;
        end else begin
          if (_T_65) begin
            out_live_in_valid_R_1_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_1_1 <= _GEN_198;
          end else begin
            if (_T_65) begin
              out_live_in_valid_R_1_1 <= 1'h0;
            end
          end
        end else begin
          if (_T_65) begin
            out_live_in_valid_R_1_1 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_1_2 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_1_2 <= _GEN_111;
        end else begin
          if (_T_66) begin
            out_live_in_valid_R_1_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_1_2 <= _GEN_199;
          end else begin
            if (_T_66) begin
              out_live_in_valid_R_1_2 <= 1'h0;
            end
          end
        end else begin
          if (_T_66) begin
            out_live_in_valid_R_1_2 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_2_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_2_0 <= _GEN_112;
        end else begin
          if (_T_67) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_2_0 <= _GEN_200;
          end else begin
            if (_T_67) begin
              out_live_in_valid_R_2_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_67) begin
            out_live_in_valid_R_2_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_3_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_3_0 <= _GEN_113;
        end else begin
          if (_T_68) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_3_0 <= _GEN_201;
          end else begin
            if (_T_68) begin
              out_live_in_valid_R_3_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_68) begin
            out_live_in_valid_R_3_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_4_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_4_0 <= _GEN_114;
        end else begin
          if (_T_69) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_4_0 <= _GEN_202;
          end else begin
            if (_T_69) begin
              out_live_in_valid_R_4_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_69) begin
            out_live_in_valid_R_4_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_5_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_5_0 <= _GEN_115;
        end else begin
          if (_T_70) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_5_0 <= _GEN_203;
          end else begin
            if (_T_70) begin
              out_live_in_valid_R_5_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_70) begin
            out_live_in_valid_R_5_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_6_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_6_0 <= _GEN_116;
        end else begin
          if (_T_71) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_6_0 <= _GEN_204;
          end else begin
            if (_T_71) begin
              out_live_in_valid_R_6_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_71) begin
            out_live_in_valid_R_6_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_7_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_7_0 <= _GEN_117;
        end else begin
          if (_T_72) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_7_0 <= _GEN_205;
          end else begin
            if (_T_72) begin
              out_live_in_valid_R_7_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_72) begin
            out_live_in_valid_R_7_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_8_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_8_0 <= _GEN_118;
        end else begin
          if (_T_73) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_8_0 <= _GEN_206;
          end else begin
            if (_T_73) begin
              out_live_in_valid_R_8_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_73) begin
            out_live_in_valid_R_8_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_9_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_9_0 <= _GEN_119;
        end else begin
          if (_T_74) begin
            out_live_in_valid_R_9_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_9_0 <= _GEN_207;
          end else begin
            if (_T_74) begin
              out_live_in_valid_R_9_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_74) begin
            out_live_in_valid_R_9_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_10_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_10_0 <= _GEN_120;
        end else begin
          if (_T_75) begin
            out_live_in_valid_R_10_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_10_0 <= _GEN_208;
          end else begin
            if (_T_75) begin
              out_live_in_valid_R_10_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_75) begin
            out_live_in_valid_R_10_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_11_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_11_0 <= _GEN_121;
        end else begin
          if (_T_76) begin
            out_live_in_valid_R_11_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_11_0 <= _GEN_209;
          end else begin
            if (_T_76) begin
              out_live_in_valid_R_11_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_76) begin
            out_live_in_valid_R_11_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_valid_R_12_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_live_in_valid_R_12_0 <= _GEN_122;
        end else begin
          if (_T_77) begin
            out_live_in_valid_R_12_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_live_in_valid_R_12_0 <= _GEN_210;
          end else begin
            if (_T_77) begin
              out_live_in_valid_R_12_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_77) begin
            out_live_in_valid_R_12_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_0_0 <= _GEN_71;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_0 <= _GEN_71;
            end
          end else begin
            out_live_in_fire_R_0_0 <= _GEN_71;
          end
        end else begin
          out_live_in_fire_R_0_0 <= _GEN_71;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_1 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_0_1 <= _GEN_73;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_1 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_1 <= _GEN_73;
            end
          end else begin
            out_live_in_fire_R_0_1 <= _GEN_73;
          end
        end else begin
          out_live_in_fire_R_0_1 <= _GEN_73;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_0_2 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_0_2 <= _GEN_75;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_0_2 <= 1'h0;
            end else begin
              out_live_in_fire_R_0_2 <= _GEN_75;
            end
          end else begin
            out_live_in_fire_R_0_2 <= _GEN_75;
          end
        end else begin
          out_live_in_fire_R_0_2 <= _GEN_75;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_1_0 <= _GEN_77;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_0 <= _GEN_77;
            end
          end else begin
            out_live_in_fire_R_1_0 <= _GEN_77;
          end
        end else begin
          out_live_in_fire_R_1_0 <= _GEN_77;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_1 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_1_1 <= _GEN_79;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_1 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_1 <= _GEN_79;
            end
          end else begin
            out_live_in_fire_R_1_1 <= _GEN_79;
          end
        end else begin
          out_live_in_fire_R_1_1 <= _GEN_79;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_1_2 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_1_2 <= _GEN_81;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_1_2 <= 1'h0;
            end else begin
              out_live_in_fire_R_1_2 <= _GEN_81;
            end
          end else begin
            out_live_in_fire_R_1_2 <= _GEN_81;
          end
        end else begin
          out_live_in_fire_R_1_2 <= _GEN_81;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_2_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_2_0 <= _GEN_83;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_2_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_2_0 <= _GEN_83;
            end
          end else begin
            out_live_in_fire_R_2_0 <= _GEN_83;
          end
        end else begin
          out_live_in_fire_R_2_0 <= _GEN_83;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_3_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_3_0 <= _GEN_85;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_3_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_3_0 <= _GEN_85;
            end
          end else begin
            out_live_in_fire_R_3_0 <= _GEN_85;
          end
        end else begin
          out_live_in_fire_R_3_0 <= _GEN_85;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_4_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_4_0 <= _GEN_87;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_4_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_4_0 <= _GEN_87;
            end
          end else begin
            out_live_in_fire_R_4_0 <= _GEN_87;
          end
        end else begin
          out_live_in_fire_R_4_0 <= _GEN_87;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_5_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_5_0 <= _GEN_89;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_5_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_5_0 <= _GEN_89;
            end
          end else begin
            out_live_in_fire_R_5_0 <= _GEN_89;
          end
        end else begin
          out_live_in_fire_R_5_0 <= _GEN_89;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_6_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_6_0 <= _GEN_91;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_6_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_6_0 <= _GEN_91;
            end
          end else begin
            out_live_in_fire_R_6_0 <= _GEN_91;
          end
        end else begin
          out_live_in_fire_R_6_0 <= _GEN_91;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_7_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_7_0 <= _GEN_93;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_7_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_7_0 <= _GEN_93;
            end
          end else begin
            out_live_in_fire_R_7_0 <= _GEN_93;
          end
        end else begin
          out_live_in_fire_R_7_0 <= _GEN_93;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_8_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_8_0 <= _GEN_95;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_8_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_8_0 <= _GEN_95;
            end
          end else begin
            out_live_in_fire_R_8_0 <= _GEN_95;
          end
        end else begin
          out_live_in_fire_R_8_0 <= _GEN_95;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_9_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_9_0 <= _GEN_97;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_9_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_9_0 <= _GEN_97;
            end
          end else begin
            out_live_in_fire_R_9_0 <= _GEN_97;
          end
        end else begin
          out_live_in_fire_R_9_0 <= _GEN_97;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_10_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_10_0 <= _GEN_99;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_10_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_10_0 <= _GEN_99;
            end
          end else begin
            out_live_in_fire_R_10_0 <= _GEN_99;
          end
        end else begin
          out_live_in_fire_R_10_0 <= _GEN_99;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_11_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_11_0 <= _GEN_101;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_11_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_11_0 <= _GEN_101;
            end
          end else begin
            out_live_in_fire_R_11_0 <= _GEN_101;
          end
        end else begin
          out_live_in_fire_R_11_0 <= _GEN_101;
        end
      end
    end
    if (reset) begin
      out_live_in_fire_R_12_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        out_live_in_fire_R_12_0 <= _GEN_103;
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              out_live_in_fire_R_12_0 <= 1'h0;
            end else begin
              out_live_in_fire_R_12_0 <= _GEN_103;
            end
          end else begin
            out_live_in_fire_R_12_0 <= _GEN_103;
          end
        end else begin
          out_live_in_fire_R_12_0 <= _GEN_103;
        end
      end
    end
    if (reset) begin
      out_carry_out_valid_R_0_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          out_carry_out_valid_R_0_0 <= _GEN_123;
        end else begin
          if (_T_78) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            out_carry_out_valid_R_0_0 <= _GEN_211;
          end else begin
            if (_T_78) begin
              out_carry_out_valid_R_0_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_78) begin
            out_carry_out_valid_R_0_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          if (enable_R_control) begin
            active_loop_start_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          active_loop_start_R_control <= _GEN_124;
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              active_loop_start_R_control <= 1'h0;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_start_R_control <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_start_valid_R <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          active_loop_start_valid_R <= _GEN_126;
        end else begin
          if (_T_58) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            active_loop_start_valid_R <= _GEN_172;
          end else begin
            if (_T_58) begin
              active_loop_start_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_58) begin
            active_loop_start_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          if (enable_R_control) begin
            active_loop_back_R_taskID <= enable_R_taskID;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              active_loop_back_R_taskID <= loop_back_R_0_taskID;
            end else begin
              if (loop_finish_R_0_control) begin
                active_loop_back_R_taskID <= 5'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_R_control <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          if (enable_R_control) begin
            active_loop_back_R_control <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            active_loop_back_R_control <= _GEN_173;
          end
        end
      end
    end
    if (reset) begin
      active_loop_back_valid_R <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          active_loop_back_valid_R <= _GEN_129;
        end else begin
          if (_T_59) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            active_loop_back_valid_R <= _GEN_175;
          end else begin
            if (_T_59) begin
              active_loop_back_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_59) begin
            active_loop_back_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_taskID <= 5'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          if (!(enable_R_control)) begin
            loop_exit_R_0_taskID <= 5'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (!(loop_back_R_0_control)) begin
              if (loop_finish_R_0_control) begin
                loop_exit_R_0_taskID <= loop_back_R_0_taskID;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_R_0_control <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          loop_exit_R_0_control <= _GEN_131;
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (!(loop_back_R_0_control)) begin
              loop_exit_R_0_control <= _GEN_167;
            end
          end
        end
      end
    end
    if (reset) begin
      loop_exit_valid_R_0 <= 1'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          if (enable_R_control) begin
            if (_T_60) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end else begin
            loop_exit_valid_R_0 <= 1'h1;
          end
        end else begin
          if (_T_60) begin
            loop_exit_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              if (_T_60) begin
                loop_exit_valid_R_0 <= 1'h0;
              end
            end else begin
              loop_exit_valid_R_0 <= _GEN_162;
            end
          end else begin
            if (_T_60) begin
              loop_exit_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          loop_exit_valid_R_0 <= _GEN_68;
        end
      end
    end
    if (reset) begin
      loop_exit_fire_R_0 <= 1'h0;
    end else begin
      loop_exit_fire_R_0 <= _GEN_69;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_79) begin
        if (_T_92) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_96) begin
          if (_T_115) begin
            if (loop_back_R_0_control) begin
              state <= 2'h1;
            end else begin
              if (loop_finish_R_0_control) begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_131) begin
            if (loop_exit_fire_R_0) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_621 & _T_123) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOOP]   Loop_1: Restarted fired @ %d\n",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 932:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_627 & _T_123) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOOP]   Loop_1: Output fired @ %d ",io_activate_loop_start_bits_taskID,value); // @[LoopBlock.scala 950:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_627 & _T_123) begin
          $fwrite(32'h80000002,"\n"); // @[LoopBlock.scala 955:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output [4:0] io_Out_5_bits_taskID,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output [4:0] io_Out_6_bits_taskID,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output [4:0] io_Out_7_bits_taskID,
  input        io_Out_8_ready,
  output       io_Out_8_valid,
  output [4:0] io_Out_8_bits_taskID,
  output       io_Out_8_bits_control,
  input        io_Out_9_ready,
  output       io_Out_9_valid,
  output [4:0] io_Out_9_bits_taskID,
  output       io_Out_9_bits_control,
  input        io_Out_10_ready,
  output       io_Out_10_valid,
  output [4:0] io_Out_10_bits_taskID,
  output       io_Out_10_bits_control,
  input        io_Out_11_ready,
  output       io_Out_11_valid,
  output [4:0] io_Out_11_bits_taskID,
  output       io_Out_11_bits_control,
  input        io_Out_12_ready,
  output       io_Out_12_valid,
  output [4:0] io_Out_12_bits_taskID,
  output       io_Out_12_bits_control,
  input        io_Out_13_ready,
  output       io_Out_13_valid,
  output [4:0] io_Out_13_bits_taskID,
  output       io_Out_13_bits_control,
  input        io_Out_14_ready,
  output       io_Out_14_valid,
  output [4:0] io_Out_14_bits_taskID,
  output       io_Out_14_bits_control,
  input        io_Out_15_ready,
  output       io_Out_15_valid,
  output [4:0] io_Out_15_bits_taskID,
  output       io_Out_15_bits_control,
  input        io_Out_16_ready,
  output       io_Out_16_valid,
  output [4:0] io_Out_16_bits_taskID,
  output       io_Out_16_bits_control,
  input        io_Out_17_ready,
  output       io_Out_17_valid,
  output [4:0] io_Out_17_bits_taskID,
  output       io_Out_17_bits_control,
  input        io_Out_18_ready,
  output       io_Out_18_valid,
  output [4:0] io_Out_18_bits_taskID,
  output       io_Out_18_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_valid_R_1; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_6;
  reg  output_valid_R_2; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_7;
  reg  output_valid_R_3; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_8;
  reg  output_valid_R_4; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_9;
  reg  output_valid_R_5; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_10;
  reg  output_valid_R_6; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_11;
  reg  output_valid_R_7; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_12;
  reg  output_valid_R_8; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_13;
  reg  output_valid_R_9; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_14;
  reg  output_valid_R_10; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_15;
  reg  output_valid_R_11; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_16;
  reg  output_valid_R_12; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_17;
  reg  output_valid_R_13; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_18;
  reg  output_valid_R_14; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_19;
  reg  output_valid_R_15; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_20;
  reg  output_valid_R_16; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_21;
  reg  output_valid_R_17; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_22;
  reg  output_valid_R_18; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_23;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_24;
  reg  output_fire_R_1; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_25;
  reg  output_fire_R_2; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_26;
  reg  output_fire_R_3; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_27;
  reg  output_fire_R_4; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_28;
  reg  output_fire_R_5; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_29;
  reg  output_fire_R_6; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_30;
  reg  output_fire_R_7; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_31;
  reg  output_fire_R_8; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_32;
  reg  output_fire_R_9; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_33;
  reg  output_fire_R_10; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_34;
  reg  output_fire_R_11; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_35;
  reg  output_fire_R_12; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_36;
  reg  output_fire_R_13; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_37;
  reg  output_fire_R_14; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_38;
  reg  output_fire_R_15; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_39;
  reg  output_fire_R_16; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_40;
  reg  output_fire_R_17; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_41;
  reg  output_fire_R_18; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_42;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BasicBlock.scala 244:28]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[BasicBlock.scala 244:28]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_10; // @[BasicBlock.scala 244:28]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_12; // @[BasicBlock.scala 244:28]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_14; // @[BasicBlock.scala 244:28]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_16; // @[BasicBlock.scala 244:28]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_18; // @[BasicBlock.scala 244:28]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[BasicBlock.scala 244:28]
  wire  _T_17; // @[Decoupled.scala 40:37]
  wire  _GEN_22; // @[BasicBlock.scala 244:28]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_24; // @[BasicBlock.scala 244:28]
  wire  _T_19; // @[Decoupled.scala 40:37]
  wire  _GEN_26; // @[BasicBlock.scala 244:28]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_28; // @[BasicBlock.scala 244:28]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_30; // @[BasicBlock.scala 244:28]
  wire  _T_22; // @[Decoupled.scala 40:37]
  wire  _GEN_32; // @[BasicBlock.scala 244:28]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _GEN_34; // @[BasicBlock.scala 244:28]
  wire  _T_24; // @[Decoupled.scala 40:37]
  wire  _GEN_36; // @[BasicBlock.scala 244:28]
  wire  _T_25; // @[Decoupled.scala 40:37]
  wire  _GEN_38; // @[BasicBlock.scala 244:28]
  wire  _T_26; // @[Decoupled.scala 40:37]
  wire  _GEN_40; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_1; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_2; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_3; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_4; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_5; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_6; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_7; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_8; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_9; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_10; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_11; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_12; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_13; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_14; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_15; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_16; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_17; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_18; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_43;
  wire  _T_69; // @[Conditional.scala 37:30]
  wire  _T_89; // @[BasicBlock.scala 309:81]
  wire  _T_90; // @[BasicBlock.scala 309:81]
  wire  _T_91; // @[BasicBlock.scala 309:81]
  wire  _T_92; // @[BasicBlock.scala 309:81]
  wire  _T_93; // @[BasicBlock.scala 309:81]
  wire  _T_94; // @[BasicBlock.scala 309:81]
  wire  _T_95; // @[BasicBlock.scala 309:81]
  wire  _T_96; // @[BasicBlock.scala 309:81]
  wire  _T_97; // @[BasicBlock.scala 309:81]
  wire  _T_98; // @[BasicBlock.scala 309:81]
  wire  _T_99; // @[BasicBlock.scala 309:81]
  wire  _T_100; // @[BasicBlock.scala 309:81]
  wire  _T_101; // @[BasicBlock.scala 309:81]
  wire  _T_102; // @[BasicBlock.scala 309:81]
  wire  _T_103; // @[BasicBlock.scala 309:81]
  wire  _T_104; // @[BasicBlock.scala 309:81]
  wire  _T_105; // @[BasicBlock.scala 309:81]
  wire  _T_106; // @[BasicBlock.scala 309:81]
  wire  _T_107; // @[BasicBlock.scala 309:81]
  wire  _T_108; // @[BasicBlock.scala 315:19]
  wire  _T_109; // @[BasicBlock.scala 315:19]
  wire  _GEN_42; // @[BasicBlock.scala 304:8]
  wire  _GEN_43; // @[BasicBlock.scala 304:8]
  wire  _GEN_44; // @[BasicBlock.scala 304:8]
  wire  _GEN_45; // @[BasicBlock.scala 304:8]
  wire  _GEN_46; // @[BasicBlock.scala 304:8]
  wire  _GEN_47; // @[BasicBlock.scala 304:8]
  wire  _GEN_48; // @[BasicBlock.scala 304:8]
  wire  _GEN_49; // @[BasicBlock.scala 304:8]
  wire  _GEN_50; // @[BasicBlock.scala 304:8]
  wire  _GEN_51; // @[BasicBlock.scala 304:8]
  wire  _GEN_52; // @[BasicBlock.scala 304:8]
  wire  _GEN_53; // @[BasicBlock.scala 304:8]
  wire  _GEN_54; // @[BasicBlock.scala 304:8]
  wire  _GEN_55; // @[BasicBlock.scala 304:8]
  wire  _GEN_56; // @[BasicBlock.scala 304:8]
  wire  _GEN_57; // @[BasicBlock.scala 304:8]
  wire  _GEN_58; // @[BasicBlock.scala 304:8]
  wire  _GEN_59; // @[BasicBlock.scala 304:8]
  wire  _GEN_60; // @[BasicBlock.scala 304:8]
  wire  _GEN_80; // @[BasicBlock.scala 304:8]
  wire  _T_113; // @[BasicBlock.scala 328:35]
  wire  _T_114; // @[BasicBlock.scala 328:35]
  wire  _T_115; // @[BasicBlock.scala 328:35]
  wire  _T_116; // @[BasicBlock.scala 328:35]
  wire  _T_117; // @[BasicBlock.scala 328:35]
  wire  _T_118; // @[BasicBlock.scala 328:35]
  wire  _T_119; // @[BasicBlock.scala 328:35]
  wire  _T_120; // @[BasicBlock.scala 328:35]
  wire  _T_121; // @[BasicBlock.scala 328:35]
  wire  _T_122; // @[BasicBlock.scala 328:35]
  wire  _T_123; // @[BasicBlock.scala 328:35]
  wire  _T_124; // @[BasicBlock.scala 328:35]
  wire  _T_125; // @[BasicBlock.scala 328:35]
  wire  _T_126; // @[BasicBlock.scala 328:35]
  wire  _T_127; // @[BasicBlock.scala 328:35]
  wire  _T_128; // @[BasicBlock.scala 328:35]
  wire  _T_129; // @[BasicBlock.scala 328:35]
  wire  _T_130; // @[BasicBlock.scala 328:35]
  wire  _GEN_188; // @[BasicBlock.scala 315:19]
  wire  _GEN_189; // @[BasicBlock.scala 315:19]
  wire  _GEN_191; // @[BasicBlock.scala 320:19]
  wire  _GEN_192; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 244:28]
  assign _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 244:28]
  assign _T_11 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_10 = _T_11 | output_fire_R_3; // @[BasicBlock.scala 244:28]
  assign _T_12 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_12 = _T_12 | output_fire_R_4; // @[BasicBlock.scala 244:28]
  assign _T_13 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_14 = _T_13 | output_fire_R_5; // @[BasicBlock.scala 244:28]
  assign _T_14 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_16 = _T_14 | output_fire_R_6; // @[BasicBlock.scala 244:28]
  assign _T_15 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_18 = _T_15 | output_fire_R_7; // @[BasicBlock.scala 244:28]
  assign _T_16 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_16 | output_fire_R_8; // @[BasicBlock.scala 244:28]
  assign _T_17 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = _T_17 | output_fire_R_9; // @[BasicBlock.scala 244:28]
  assign _T_18 = io_Out_10_ready & io_Out_10_valid; // @[Decoupled.scala 40:37]
  assign _GEN_24 = _T_18 | output_fire_R_10; // @[BasicBlock.scala 244:28]
  assign _T_19 = io_Out_11_ready & io_Out_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_26 = _T_19 | output_fire_R_11; // @[BasicBlock.scala 244:28]
  assign _T_20 = io_Out_12_ready & io_Out_12_valid; // @[Decoupled.scala 40:37]
  assign _GEN_28 = _T_20 | output_fire_R_12; // @[BasicBlock.scala 244:28]
  assign _T_21 = io_Out_13_ready & io_Out_13_valid; // @[Decoupled.scala 40:37]
  assign _GEN_30 = _T_21 | output_fire_R_13; // @[BasicBlock.scala 244:28]
  assign _T_22 = io_Out_14_ready & io_Out_14_valid; // @[Decoupled.scala 40:37]
  assign _GEN_32 = _T_22 | output_fire_R_14; // @[BasicBlock.scala 244:28]
  assign _T_23 = io_Out_15_ready & io_Out_15_valid; // @[Decoupled.scala 40:37]
  assign _GEN_34 = _T_23 | output_fire_R_15; // @[BasicBlock.scala 244:28]
  assign _T_24 = io_Out_16_ready & io_Out_16_valid; // @[Decoupled.scala 40:37]
  assign _GEN_36 = _T_24 | output_fire_R_16; // @[BasicBlock.scala 244:28]
  assign _T_25 = io_Out_17_ready & io_Out_17_valid; // @[Decoupled.scala 40:37]
  assign _GEN_38 = _T_25 | output_fire_R_17; // @[BasicBlock.scala 244:28]
  assign _T_26 = io_Out_18_ready & io_Out_18_valid; // @[Decoupled.scala 40:37]
  assign _GEN_40 = _T_26 | output_fire_R_18; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_3 = output_fire_R_3 | _T_11; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_4 = output_fire_R_4 | _T_12; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_5 = output_fire_R_5 | _T_13; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_6 = output_fire_R_6 | _T_14; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_7 = output_fire_R_7 | _T_15; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_8 = output_fire_R_8 | _T_16; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_9 = output_fire_R_9 | _T_17; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_10 = output_fire_R_10 | _T_18; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_11 = output_fire_R_11 | _T_19; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_12 = output_fire_R_12 | _T_20; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_13 = output_fire_R_13 | _T_21; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_14 = output_fire_R_14 | _T_22; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_15 = output_fire_R_15 | _T_23; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_16 = output_fire_R_16 | _T_24; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_17 = output_fire_R_17 | _T_25; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_18 = output_fire_R_18 | _T_26; // @[BasicBlock.scala 256:85]
  assign _T_69 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_89 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_90 = _T_9 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_91 = _T_10 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_92 = _T_11 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_93 = _T_12 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_94 = _T_13 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_95 = _T_14 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_96 = _T_15 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_97 = _T_16 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_98 = _T_17 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_99 = _T_18 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_100 = _T_19 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_101 = _T_20 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_102 = _T_21 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_103 = _T_22 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_104 = _T_23 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_105 = _T_24 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_106 = _T_25 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_107 = _T_26 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_108 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_109 = _T_108 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_42 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_43 = _GEN_3 | output_valid_R_1; // @[BasicBlock.scala 304:8]
  assign _GEN_44 = _GEN_3 | output_valid_R_2; // @[BasicBlock.scala 304:8]
  assign _GEN_45 = _GEN_3 | output_valid_R_3; // @[BasicBlock.scala 304:8]
  assign _GEN_46 = _GEN_3 | output_valid_R_4; // @[BasicBlock.scala 304:8]
  assign _GEN_47 = _GEN_3 | output_valid_R_5; // @[BasicBlock.scala 304:8]
  assign _GEN_48 = _GEN_3 | output_valid_R_6; // @[BasicBlock.scala 304:8]
  assign _GEN_49 = _GEN_3 | output_valid_R_7; // @[BasicBlock.scala 304:8]
  assign _GEN_50 = _GEN_3 | output_valid_R_8; // @[BasicBlock.scala 304:8]
  assign _GEN_51 = _GEN_3 | output_valid_R_9; // @[BasicBlock.scala 304:8]
  assign _GEN_52 = _GEN_3 | output_valid_R_10; // @[BasicBlock.scala 304:8]
  assign _GEN_53 = _GEN_3 | output_valid_R_11; // @[BasicBlock.scala 304:8]
  assign _GEN_54 = _GEN_3 | output_valid_R_12; // @[BasicBlock.scala 304:8]
  assign _GEN_55 = _GEN_3 | output_valid_R_13; // @[BasicBlock.scala 304:8]
  assign _GEN_56 = _GEN_3 | output_valid_R_14; // @[BasicBlock.scala 304:8]
  assign _GEN_57 = _GEN_3 | output_valid_R_15; // @[BasicBlock.scala 304:8]
  assign _GEN_58 = _GEN_3 | output_valid_R_16; // @[BasicBlock.scala 304:8]
  assign _GEN_59 = _GEN_3 | output_valid_R_17; // @[BasicBlock.scala 304:8]
  assign _GEN_60 = _GEN_3 | output_valid_R_18; // @[BasicBlock.scala 304:8]
  assign _GEN_80 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign _T_113 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 328:35]
  assign _T_114 = _T_113 & out_fire_mask_2; // @[BasicBlock.scala 328:35]
  assign _T_115 = _T_114 & out_fire_mask_3; // @[BasicBlock.scala 328:35]
  assign _T_116 = _T_115 & out_fire_mask_4; // @[BasicBlock.scala 328:35]
  assign _T_117 = _T_116 & out_fire_mask_5; // @[BasicBlock.scala 328:35]
  assign _T_118 = _T_117 & out_fire_mask_6; // @[BasicBlock.scala 328:35]
  assign _T_119 = _T_118 & out_fire_mask_7; // @[BasicBlock.scala 328:35]
  assign _T_120 = _T_119 & out_fire_mask_8; // @[BasicBlock.scala 328:35]
  assign _T_121 = _T_120 & out_fire_mask_9; // @[BasicBlock.scala 328:35]
  assign _T_122 = _T_121 & out_fire_mask_10; // @[BasicBlock.scala 328:35]
  assign _T_123 = _T_122 & out_fire_mask_11; // @[BasicBlock.scala 328:35]
  assign _T_124 = _T_123 & out_fire_mask_12; // @[BasicBlock.scala 328:35]
  assign _T_125 = _T_124 & out_fire_mask_13; // @[BasicBlock.scala 328:35]
  assign _T_126 = _T_125 & out_fire_mask_14; // @[BasicBlock.scala 328:35]
  assign _T_127 = _T_126 & out_fire_mask_15; // @[BasicBlock.scala 328:35]
  assign _T_128 = _T_127 & out_fire_mask_16; // @[BasicBlock.scala 328:35]
  assign _T_129 = _T_128 & out_fire_mask_17; // @[BasicBlock.scala 328:35]
  assign _T_130 = _T_129 & out_fire_mask_18; // @[BasicBlock.scala 328:35]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_69 ? _GEN_42 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_1_valid = _T_69 ? _GEN_43 : output_valid_R_1; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_2_valid = _T_69 ? _GEN_44 : output_valid_R_2; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_3_valid = _T_69 ? _GEN_45 : output_valid_R_3; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_3_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_4_valid = _T_69 ? _GEN_46 : output_valid_R_4; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_4_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_5_valid = _T_69 ? _GEN_47 : output_valid_R_5; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_5_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_6_valid = _T_69 ? _GEN_48 : output_valid_R_6; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_6_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_7_valid = _T_69 ? _GEN_49 : output_valid_R_7; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_7_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_8_valid = _T_69 ? _GEN_50 : output_valid_R_8; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_8_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_8_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_9_valid = _T_69 ? _GEN_51 : output_valid_R_9; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_9_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_9_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_10_valid = _T_69 ? _GEN_52 : output_valid_R_10; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_10_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_10_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_11_valid = _T_69 ? _GEN_53 : output_valid_R_11; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_11_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_11_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_12_valid = _T_69 ? _GEN_54 : output_valid_R_12; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_12_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_12_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_13_valid = _T_69 ? _GEN_55 : output_valid_R_13; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_13_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_13_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_14_valid = _T_69 ? _GEN_56 : output_valid_R_14; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_14_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_14_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_15_valid = _T_69 ? _GEN_57 : output_valid_R_15; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_15_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_15_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_16_valid = _T_69 ? _GEN_58 : output_valid_R_16; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_16_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_16_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_17_valid = _T_69 ? _GEN_59 : output_valid_R_17; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_17_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_17_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_18_valid = _T_69 ? _GEN_60 : output_valid_R_18; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_18_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_18_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_188 = _T_69 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_189 = _GEN_188 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_191 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_192 = _GEN_188 & _GEN_191; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_4 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_valid_R_5 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_valid_R_6 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_valid_R_7 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  output_valid_R_8 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  output_valid_R_9 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  output_valid_R_10 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  output_valid_R_11 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  output_valid_R_12 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  output_valid_R_13 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  output_valid_R_14 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  output_valid_R_15 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  output_valid_R_16 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  output_valid_R_17 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  output_valid_R_18 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  output_fire_R_4 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  output_fire_R_5 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  output_fire_R_6 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  output_fire_R_7 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  output_fire_R_8 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  output_fire_R_9 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  output_fire_R_10 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  output_fire_R_11 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  output_fire_R_12 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  output_fire_R_13 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  output_fire_R_14 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  output_fire_R_15 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  output_fire_R_16 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  output_fire_R_17 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  output_fire_R_18 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  state = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_69) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_130) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_130) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_69) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_130) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_89;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_1 <= _T_90;
        end else begin
          if (_T_9) begin
            output_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_9) begin
          output_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_2 <= _T_91;
        end else begin
          if (_T_10) begin
            output_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_10) begin
          output_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_3 <= _T_92;
        end else begin
          if (_T_11) begin
            output_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_11) begin
          output_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_4 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_4 <= _T_93;
        end else begin
          if (_T_12) begin
            output_valid_R_4 <= 1'h0;
          end
        end
      end else begin
        if (_T_12) begin
          output_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_5 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_5 <= _T_94;
        end else begin
          if (_T_13) begin
            output_valid_R_5 <= 1'h0;
          end
        end
      end else begin
        if (_T_13) begin
          output_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_6 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_6 <= _T_95;
        end else begin
          if (_T_14) begin
            output_valid_R_6 <= 1'h0;
          end
        end
      end else begin
        if (_T_14) begin
          output_valid_R_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_7 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_7 <= _T_96;
        end else begin
          if (_T_15) begin
            output_valid_R_7 <= 1'h0;
          end
        end
      end else begin
        if (_T_15) begin
          output_valid_R_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_8 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_8 <= _T_97;
        end else begin
          if (_T_16) begin
            output_valid_R_8 <= 1'h0;
          end
        end
      end else begin
        if (_T_16) begin
          output_valid_R_8 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_9 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_9 <= _T_98;
        end else begin
          if (_T_17) begin
            output_valid_R_9 <= 1'h0;
          end
        end
      end else begin
        if (_T_17) begin
          output_valid_R_9 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_10 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_10 <= _T_99;
        end else begin
          if (_T_18) begin
            output_valid_R_10 <= 1'h0;
          end
        end
      end else begin
        if (_T_18) begin
          output_valid_R_10 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_11 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_11 <= _T_100;
        end else begin
          if (_T_19) begin
            output_valid_R_11 <= 1'h0;
          end
        end
      end else begin
        if (_T_19) begin
          output_valid_R_11 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_12 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_12 <= _T_101;
        end else begin
          if (_T_20) begin
            output_valid_R_12 <= 1'h0;
          end
        end
      end else begin
        if (_T_20) begin
          output_valid_R_12 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_13 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_13 <= _T_102;
        end else begin
          if (_T_21) begin
            output_valid_R_13 <= 1'h0;
          end
        end
      end else begin
        if (_T_21) begin
          output_valid_R_13 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_14 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_14 <= _T_103;
        end else begin
          if (_T_22) begin
            output_valid_R_14 <= 1'h0;
          end
        end
      end else begin
        if (_T_22) begin
          output_valid_R_14 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_15 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_15 <= _T_104;
        end else begin
          if (_T_23) begin
            output_valid_R_15 <= 1'h0;
          end
        end
      end else begin
        if (_T_23) begin
          output_valid_R_15 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_16 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_16 <= _T_105;
        end else begin
          if (_T_24) begin
            output_valid_R_16 <= 1'h0;
          end
        end
      end else begin
        if (_T_24) begin
          output_valid_R_16 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_17 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_17 <= _T_106;
        end else begin
          if (_T_25) begin
            output_valid_R_17 <= 1'h0;
          end
        end
      end else begin
        if (_T_25) begin
          output_valid_R_17 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_18 <= 1'h0;
    end else begin
      if (_T_69) begin
        if (_GEN_3) begin
          output_valid_R_18 <= _T_107;
        end else begin
          if (_T_26) begin
            output_valid_R_18 <= 1'h0;
          end
        end
      end else begin
        if (_T_26) begin
          output_valid_R_18 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_1 <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_1 <= 1'h0;
          end else begin
            output_fire_R_1 <= _GEN_6;
          end
        end else begin
          output_fire_R_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_2 <= _GEN_8;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_2 <= 1'h0;
          end else begin
            output_fire_R_2 <= _GEN_8;
          end
        end else begin
          output_fire_R_2 <= _GEN_8;
        end
      end
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_3 <= _GEN_10;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_3 <= 1'h0;
          end else begin
            output_fire_R_3 <= _GEN_10;
          end
        end else begin
          output_fire_R_3 <= _GEN_10;
        end
      end
    end
    if (reset) begin
      output_fire_R_4 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_4 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_4 <= 1'h0;
          end else begin
            output_fire_R_4 <= _GEN_12;
          end
        end else begin
          output_fire_R_4 <= _GEN_12;
        end
      end
    end
    if (reset) begin
      output_fire_R_5 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_5 <= _GEN_14;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_5 <= 1'h0;
          end else begin
            output_fire_R_5 <= _GEN_14;
          end
        end else begin
          output_fire_R_5 <= _GEN_14;
        end
      end
    end
    if (reset) begin
      output_fire_R_6 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_6 <= _GEN_16;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_6 <= 1'h0;
          end else begin
            output_fire_R_6 <= _GEN_16;
          end
        end else begin
          output_fire_R_6 <= _GEN_16;
        end
      end
    end
    if (reset) begin
      output_fire_R_7 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_7 <= _GEN_18;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_7 <= 1'h0;
          end else begin
            output_fire_R_7 <= _GEN_18;
          end
        end else begin
          output_fire_R_7 <= _GEN_18;
        end
      end
    end
    if (reset) begin
      output_fire_R_8 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_8 <= _GEN_20;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_8 <= 1'h0;
          end else begin
            output_fire_R_8 <= _GEN_20;
          end
        end else begin
          output_fire_R_8 <= _GEN_20;
        end
      end
    end
    if (reset) begin
      output_fire_R_9 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_9 <= _GEN_22;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_9 <= 1'h0;
          end else begin
            output_fire_R_9 <= _GEN_22;
          end
        end else begin
          output_fire_R_9 <= _GEN_22;
        end
      end
    end
    if (reset) begin
      output_fire_R_10 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_10 <= _GEN_24;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_10 <= 1'h0;
          end else begin
            output_fire_R_10 <= _GEN_24;
          end
        end else begin
          output_fire_R_10 <= _GEN_24;
        end
      end
    end
    if (reset) begin
      output_fire_R_11 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_11 <= _GEN_26;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_11 <= 1'h0;
          end else begin
            output_fire_R_11 <= _GEN_26;
          end
        end else begin
          output_fire_R_11 <= _GEN_26;
        end
      end
    end
    if (reset) begin
      output_fire_R_12 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_12 <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_12 <= 1'h0;
          end else begin
            output_fire_R_12 <= _GEN_28;
          end
        end else begin
          output_fire_R_12 <= _GEN_28;
        end
      end
    end
    if (reset) begin
      output_fire_R_13 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_13 <= _GEN_30;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_13 <= 1'h0;
          end else begin
            output_fire_R_13 <= _GEN_30;
          end
        end else begin
          output_fire_R_13 <= _GEN_30;
        end
      end
    end
    if (reset) begin
      output_fire_R_14 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_14 <= _GEN_32;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_14 <= 1'h0;
          end else begin
            output_fire_R_14 <= _GEN_32;
          end
        end else begin
          output_fire_R_14 <= _GEN_32;
        end
      end
    end
    if (reset) begin
      output_fire_R_15 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_15 <= _GEN_34;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_15 <= 1'h0;
          end else begin
            output_fire_R_15 <= _GEN_34;
          end
        end else begin
          output_fire_R_15 <= _GEN_34;
        end
      end
    end
    if (reset) begin
      output_fire_R_16 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_16 <= _GEN_36;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_16 <= 1'h0;
          end else begin
            output_fire_R_16 <= _GEN_36;
          end
        end else begin
          output_fire_R_16 <= _GEN_36;
        end
      end
    end
    if (reset) begin
      output_fire_R_17 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_17 <= _GEN_38;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_17 <= 1'h0;
          end else begin
            output_fire_R_17 <= _GEN_38;
          end
        end else begin
          output_fire_R_17 <= _GEN_38;
        end
      end
    end
    if (reset) begin
      output_fire_R_18 <= 1'h0;
    end else begin
      if (_T_69) begin
        output_fire_R_18 <= _GEN_40;
      end else begin
        if (state) begin
          if (_T_130) begin
            output_fire_R_18 <= 1'h0;
          end else begin
            output_fire_R_18 <= _GEN_40;
          end
        end else begin
          output_fire_R_18 <= _GEN_40;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_69) begin
        state <= _GEN_80;
      end else begin
        if (state) begin
          if (_T_130) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_189 & _T_109) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [BB]   bb_entry0: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_192 & _T_109) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [BB]   bb_entry0: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_1(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_6;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_7;
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_17; // @[BasicBlock.scala 309:81]
  wire  _T_18; // @[BasicBlock.scala 315:19]
  wire  _T_19; // @[BasicBlock.scala 315:19]
  wire  _GEN_6; // @[BasicBlock.scala 304:8]
  wire  _GEN_8; // @[BasicBlock.scala 304:8]
  wire  _GEN_26; // @[BasicBlock.scala 315:19]
  wire  _GEN_27; // @[BasicBlock.scala 315:19]
  wire  _GEN_29; // @[BasicBlock.scala 320:19]
  wire  _GEN_30; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_18 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_19 = _T_18 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_6 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_8 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_15 ? _GEN_6 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_0_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_26 = _T_15 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_27 = _GEN_26 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_29 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_17;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_8;
      end else begin
        if (state) begin
          if (out_fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [BB]   bb_for_cond_cleanup1: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [BB]   bb_for_cond_cleanup1: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output       io_Out_5_bits_control,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output [4:0] io_Out_6_bits_taskID,
  output       io_Out_6_bits_control,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output [4:0] io_Out_7_bits_taskID,
  output       io_Out_7_bits_control,
  input        io_Out_8_ready,
  output       io_Out_8_valid,
  output [4:0] io_Out_8_bits_taskID,
  output       io_Out_8_bits_control,
  input        io_Out_9_ready,
  output       io_Out_9_valid,
  output [4:0] io_Out_9_bits_taskID,
  output       io_Out_9_bits_control,
  input        io_Out_10_ready,
  output       io_Out_10_valid,
  output [4:0] io_Out_10_bits_taskID,
  output       io_Out_10_bits_control,
  input        io_Out_11_ready,
  output       io_Out_11_valid,
  output [4:0] io_Out_11_bits_taskID,
  output       io_Out_11_bits_control,
  input        io_Out_12_ready,
  output       io_Out_12_valid,
  output [4:0] io_Out_12_bits_taskID,
  output       io_Out_12_bits_control,
  input        io_Out_13_ready,
  output       io_Out_13_valid,
  output [4:0] io_Out_13_bits_taskID,
  output       io_Out_13_bits_control,
  input        io_Out_14_ready,
  output       io_Out_14_valid,
  output [4:0] io_Out_14_bits_taskID,
  output       io_Out_14_bits_control,
  input        io_Out_15_ready,
  output       io_Out_15_valid,
  output [4:0] io_Out_15_bits_taskID,
  output       io_Out_15_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_4;
  reg  out_ready_R_5; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_5;
  reg  out_ready_R_6; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_6;
  reg  out_ready_R_7; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_7;
  reg  out_ready_R_8; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_8;
  reg  out_ready_R_9; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_9;
  reg  out_ready_R_10; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_10;
  reg  out_ready_R_11; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_11;
  reg  out_ready_R_12; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_12;
  reg  out_ready_R_13; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_13;
  reg  out_ready_R_14; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_14;
  reg  out_ready_R_15; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_15;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_16;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_17;
  reg  out_valid_R_2; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_18;
  reg  out_valid_R_3; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_19;
  reg  out_valid_R_4; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_20;
  reg  out_valid_R_5; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_21;
  reg  out_valid_R_6; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_22;
  reg  out_valid_R_7; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_23;
  reg  out_valid_R_8; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_24;
  reg  out_valid_R_9; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_25;
  reg  out_valid_R_10; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_26;
  reg  out_valid_R_11; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_27;
  reg  out_valid_R_12; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_28;
  reg  out_valid_R_13; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_29;
  reg  out_valid_R_14; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_30;
  reg  out_valid_R_15; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_31;
  reg  mask_valid_R_0; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_32;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 716:29]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[HandShaking.scala 716:29]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[HandShaking.scala 716:29]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[HandShaking.scala 716:29]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[HandShaking.scala 716:29]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[HandShaking.scala 716:29]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[HandShaking.scala 716:29]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[HandShaking.scala 716:29]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[HandShaking.scala 716:29]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_23; // @[HandShaking.scala 716:29]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[HandShaking.scala 716:29]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_27; // @[HandShaking.scala 716:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[HandShaking.scala 716:29]
  wire  _T_17; // @[Decoupled.scala 40:37]
  wire  _GEN_31; // @[HandShaking.scala 716:29]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[HandShaking.scala 727:32]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_33;
  wire [14:0] _T_21; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_34;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_35;
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_36;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_37;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_38;
  reg  predicate_control_R_1; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_39;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_40;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_41;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_42;
  wire  predicate; // @[BasicBlock.scala 75:58]
  wire [4:0] predicate_task; // @[BasicBlock.scala 76:62]
  wire  _T_26; // @[Decoupled.scala 40:37]
  wire  _T_27; // @[Decoupled.scala 40:37]
  wire  _T_28; // @[BasicBlock.scala 78:91]
  wire  _T_29; // @[BasicBlock.scala 78:91]
  wire  start; // @[BasicBlock.scala 78:107]
  wire [1:0] _T_34; // @[BasicBlock.scala 102:52]
  wire  _T_35; // @[Conditional.scala 37:30]
  wire  _GEN_43; // @[BasicBlock.scala 112:19]
  wire  _GEN_44; // @[BasicBlock.scala 112:19]
  wire  _GEN_45; // @[BasicBlock.scala 112:19]
  wire  _GEN_46; // @[BasicBlock.scala 112:19]
  wire  _GEN_47; // @[BasicBlock.scala 112:19]
  wire  _GEN_48; // @[BasicBlock.scala 112:19]
  wire  _GEN_49; // @[BasicBlock.scala 112:19]
  wire  _GEN_50; // @[BasicBlock.scala 112:19]
  wire  _GEN_51; // @[BasicBlock.scala 112:19]
  wire  _GEN_52; // @[BasicBlock.scala 112:19]
  wire  _GEN_53; // @[BasicBlock.scala 112:19]
  wire  _GEN_54; // @[BasicBlock.scala 112:19]
  wire  _GEN_55; // @[BasicBlock.scala 112:19]
  wire  _GEN_56; // @[BasicBlock.scala 112:19]
  wire  _GEN_57; // @[BasicBlock.scala 112:19]
  wire  _GEN_58; // @[BasicBlock.scala 112:19]
  wire  _GEN_59; // @[BasicBlock.scala 112:19]
  wire  _GEN_60; // @[BasicBlock.scala 112:19]
  wire [7:0] _T_44; // @[HandShaking.scala 741:17]
  wire [15:0] _T_52; // @[HandShaking.scala 741:17]
  wire  _T_53; // @[HandShaking.scala 741:24]
  wire  _T_56; // @[BasicBlock.scala 126:19]
  wire  _T_57; // @[BasicBlock.scala 126:19]
  wire  _GEN_138; // @[BasicBlock.scala 126:19]
  wire  _GEN_139; // @[BasicBlock.scala 126:19]
  wire  _GEN_140; // @[BasicBlock.scala 126:19]
  wire  _GEN_141; // @[BasicBlock.scala 126:19]
  wire  _GEN_145; // @[BasicBlock.scala 132:19]
  wire  _GEN_146; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 716:29]
  assign _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 716:29]
  assign _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 716:29]
  assign _T_7 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_7 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 716:29]
  assign _T_8 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_8 ? 1'h0 : out_valid_R_6; // @[HandShaking.scala 716:29]
  assign _T_9 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_9 ? 1'h0 : out_valid_R_7; // @[HandShaking.scala 716:29]
  assign _T_10 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_10 ? 1'h0 : out_valid_R_8; // @[HandShaking.scala 716:29]
  assign _T_11 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_11 ? 1'h0 : out_valid_R_9; // @[HandShaking.scala 716:29]
  assign _T_12 = io_Out_10_ready & io_Out_10_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_12 ? 1'h0 : out_valid_R_10; // @[HandShaking.scala 716:29]
  assign _T_13 = io_Out_11_ready & io_Out_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_23 = _T_13 ? 1'h0 : out_valid_R_11; // @[HandShaking.scala 716:29]
  assign _T_14 = io_Out_12_ready & io_Out_12_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_14 ? 1'h0 : out_valid_R_12; // @[HandShaking.scala 716:29]
  assign _T_15 = io_Out_13_ready & io_Out_13_valid; // @[Decoupled.scala 40:37]
  assign _GEN_27 = _T_15 ? 1'h0 : out_valid_R_13; // @[HandShaking.scala 716:29]
  assign _T_16 = io_Out_14_ready & io_Out_14_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_16 ? 1'h0 : out_valid_R_14; // @[HandShaking.scala 716:29]
  assign _T_17 = io_Out_15_ready & io_Out_15_valid; // @[Decoupled.scala 40:37]
  assign _GEN_31 = _T_17 ? 1'h0 : out_valid_R_15; // @[HandShaking.scala 716:29]
  assign _T_18 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_18 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 727:32]
  assign _T_21 = value + 15'h1; // @[Counter.scala 38:22]
  assign predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 75:58]
  assign predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 76:62]
  assign _T_26 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _T_27 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _T_28 = _T_26 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_29 = _T_27 | predicate_valid_R_1; // @[BasicBlock.scala 78:91]
  assign start = _T_28 & _T_29; // @[BasicBlock.scala 78:107]
  assign _T_34 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:52]
  assign _T_35 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_43 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_44 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_45 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_46 = start | _GEN_7; // @[BasicBlock.scala 112:19]
  assign _GEN_47 = start | _GEN_9; // @[BasicBlock.scala 112:19]
  assign _GEN_48 = start | _GEN_11; // @[BasicBlock.scala 112:19]
  assign _GEN_49 = start | _GEN_13; // @[BasicBlock.scala 112:19]
  assign _GEN_50 = start | _GEN_15; // @[BasicBlock.scala 112:19]
  assign _GEN_51 = start | _GEN_17; // @[BasicBlock.scala 112:19]
  assign _GEN_52 = start | _GEN_19; // @[BasicBlock.scala 112:19]
  assign _GEN_53 = start | _GEN_21; // @[BasicBlock.scala 112:19]
  assign _GEN_54 = start | _GEN_23; // @[BasicBlock.scala 112:19]
  assign _GEN_55 = start | _GEN_25; // @[BasicBlock.scala 112:19]
  assign _GEN_56 = start | _GEN_27; // @[BasicBlock.scala 112:19]
  assign _GEN_57 = start | _GEN_29; // @[BasicBlock.scala 112:19]
  assign _GEN_58 = start | _GEN_31; // @[BasicBlock.scala 112:19]
  assign _GEN_59 = start | _GEN_33; // @[BasicBlock.scala 112:19]
  assign _GEN_60 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_44 = {out_ready_R_7,out_ready_R_6,out_ready_R_5,out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_52 = {out_ready_R_15,out_ready_R_14,out_ready_R_13,out_ready_R_12,out_ready_R_11,out_ready_R_10,out_ready_R_9,out_ready_R_8,_T_44}; // @[HandShaking.scala 741:17]
  assign _T_53 = _T_52 == 16'hffff; // @[HandShaking.scala 741:24]
  assign _T_56 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_57 = _T_56 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 726:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 715:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 715:21]
  assign io_Out_3_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 715:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 715:21]
  assign io_Out_5_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 715:21]
  assign io_Out_6_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_6_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 715:21]
  assign io_Out_7_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_7_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_8_valid = out_valid_R_8; // @[HandShaking.scala 715:21]
  assign io_Out_8_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_8_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_9_valid = out_valid_R_9; // @[HandShaking.scala 715:21]
  assign io_Out_9_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_9_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_10_valid = out_valid_R_10; // @[HandShaking.scala 715:21]
  assign io_Out_10_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_10_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_11_valid = out_valid_R_11; // @[HandShaking.scala 715:21]
  assign io_Out_11_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_11_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_12_valid = out_valid_R_12; // @[HandShaking.scala 715:21]
  assign io_Out_12_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_12_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_13_valid = out_valid_R_13; // @[HandShaking.scala 715:21]
  assign io_Out_13_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_13_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_14_valid = out_valid_R_14; // @[HandShaking.scala 715:21]
  assign io_Out_14_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_14_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_15_valid = out_valid_R_15; // @[HandShaking.scala 715:21]
  assign io_Out_15_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_15_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 86:29]
  assign _GEN_138 = _T_35 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_139 = _GEN_138 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_140 = _GEN_139 & _T_53; // @[BasicBlock.scala 126:19]
  assign _GEN_141 = _GEN_140 & predicate; // @[BasicBlock.scala 126:19]
  assign _GEN_145 = predicate == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_146 = _GEN_140 & _GEN_145; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_ready_R_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_ready_R_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_ready_R_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_ready_R_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_ready_R_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_ready_R_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  out_ready_R_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_ready_R_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  out_valid_R_8 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  out_valid_R_9 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  out_valid_R_10 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_valid_R_11 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_valid_R_12 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_valid_R_13 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_valid_R_14 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  out_valid_R_15 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  value = _RAND_33[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_36[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  state = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_4) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_5) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_6) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_6) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_6) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_7) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_7) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_7) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_8) begin
          out_ready_R_6 <= io_Out_6_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_6 <= 1'h0;
          end else begin
            if (_T_8) begin
              out_ready_R_6 <= io_Out_6_ready;
            end
          end
        end else begin
          if (_T_8) begin
            out_ready_R_6 <= io_Out_6_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_9) begin
          out_ready_R_7 <= io_Out_7_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_7 <= 1'h0;
          end else begin
            if (_T_9) begin
              out_ready_R_7 <= io_Out_7_ready;
            end
          end
        end else begin
          if (_T_9) begin
            out_ready_R_7 <= io_Out_7_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_8 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_10) begin
          out_ready_R_8 <= io_Out_8_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_8 <= 1'h0;
          end else begin
            if (_T_10) begin
              out_ready_R_8 <= io_Out_8_ready;
            end
          end
        end else begin
          if (_T_10) begin
            out_ready_R_8 <= io_Out_8_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_9 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_11) begin
          out_ready_R_9 <= io_Out_9_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_9 <= 1'h0;
          end else begin
            if (_T_11) begin
              out_ready_R_9 <= io_Out_9_ready;
            end
          end
        end else begin
          if (_T_11) begin
            out_ready_R_9 <= io_Out_9_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_10 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_12) begin
          out_ready_R_10 <= io_Out_10_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_10 <= 1'h0;
          end else begin
            if (_T_12) begin
              out_ready_R_10 <= io_Out_10_ready;
            end
          end
        end else begin
          if (_T_12) begin
            out_ready_R_10 <= io_Out_10_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_11 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_13) begin
          out_ready_R_11 <= io_Out_11_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_11 <= 1'h0;
          end else begin
            if (_T_13) begin
              out_ready_R_11 <= io_Out_11_ready;
            end
          end
        end else begin
          if (_T_13) begin
            out_ready_R_11 <= io_Out_11_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_12 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_14) begin
          out_ready_R_12 <= io_Out_12_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_12 <= 1'h0;
          end else begin
            if (_T_14) begin
              out_ready_R_12 <= io_Out_12_ready;
            end
          end
        end else begin
          if (_T_14) begin
            out_ready_R_12 <= io_Out_12_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_13 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_15) begin
          out_ready_R_13 <= io_Out_13_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_13 <= 1'h0;
          end else begin
            if (_T_15) begin
              out_ready_R_13 <= io_Out_13_ready;
            end
          end
        end else begin
          if (_T_15) begin
            out_ready_R_13 <= io_Out_13_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_14 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_16) begin
          out_ready_R_14 <= io_Out_14_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_14 <= 1'h0;
          end else begin
            if (_T_16) begin
              out_ready_R_14 <= io_Out_14_ready;
            end
          end
        end else begin
          if (_T_16) begin
            out_ready_R_14 <= io_Out_14_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_15 <= 1'h0;
    end else begin
      if (_T_35) begin
        if (_T_17) begin
          out_ready_R_15 <= io_Out_15_ready;
        end
      end else begin
        if (state) begin
          if (_T_53) begin
            out_ready_R_15 <= 1'h0;
          end else begin
            if (_T_17) begin
              out_ready_R_15 <= io_Out_15_ready;
            end
          end
        end else begin
          if (_T_17) begin
            out_ready_R_15 <= io_Out_15_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_0 <= _GEN_43;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_1 <= _GEN_44;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_2 <= _GEN_45;
      end else begin
        if (_T_4) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_3 <= _GEN_46;
      end else begin
        if (_T_5) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_4 <= _GEN_47;
      end else begin
        if (_T_6) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_5 <= _GEN_48;
      end else begin
        if (_T_7) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_6 <= _GEN_49;
      end else begin
        if (_T_8) begin
          out_valid_R_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_7 <= _GEN_50;
      end else begin
        if (_T_9) begin
          out_valid_R_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_8 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_8 <= _GEN_51;
      end else begin
        if (_T_10) begin
          out_valid_R_8 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_9 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_9 <= _GEN_52;
      end else begin
        if (_T_11) begin
          out_valid_R_9 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_10 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_10 <= _GEN_53;
      end else begin
        if (_T_12) begin
          out_valid_R_10 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_11 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_11 <= _GEN_54;
      end else begin
        if (_T_13) begin
          out_valid_R_11 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_12 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_12 <= _GEN_55;
      end else begin
        if (_T_14) begin
          out_valid_R_12 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_13 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_13 <= _GEN_56;
      end else begin
        if (_T_15) begin
          out_valid_R_13 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_14 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_14 <= _GEN_57;
      end else begin
        if (_T_16) begin
          out_valid_R_14 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_15 <= 1'h0;
    end else begin
      if (_T_35) begin
        out_valid_R_15 <= _GEN_58;
      end else begin
        if (_T_17) begin
          out_valid_R_15 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_35) begin
        mask_valid_R_0 <= _GEN_59;
      end else begin
        if (_T_18) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_21;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_26) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_26) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_27) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_26) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_35) begin
        predicate_valid_R_0 <= _T_28;
      end else begin
        if (state) begin
          if (_T_53) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= _T_28;
          end
        end else begin
          predicate_valid_R_0 <= _T_28;
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_35) begin
        predicate_valid_R_1 <= _T_29;
      end else begin
        if (state) begin
          if (_T_53) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            predicate_valid_R_1 <= _T_29;
          end
        end else begin
          predicate_valid_R_1 <= _T_29;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_35) begin
        state <= _GEN_60;
      end else begin
        if (state) begin
          if (_T_53) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_141 & _T_57) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [BB]   bb_for_body2: Output fired @ %d, Mask: %d\n",predicate_task,value,_T_34); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_146 & _T_57) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] bb_for_body2: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNoMaskFastNode_2(
  input        clock,
  input        reset,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  output       io_Out_2_bits_control,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  output       io_Out_3_bits_control,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  output       io_Out_4_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] in_data_R_0_taskID; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_1;
  reg  in_data_R_0_control; // @[BasicBlock.scala 222:46]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_0; // @[BasicBlock.scala 223:52]
  reg [31:0] _RAND_3;
  reg [4:0] output_R_taskID; // @[BasicBlock.scala 225:25]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_5;
  reg  output_valid_R_1; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_6;
  reg  output_valid_R_2; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_7;
  reg  output_valid_R_3; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_8;
  reg  output_valid_R_4; // @[BasicBlock.scala 226:49]
  reg [31:0] _RAND_9;
  reg  output_fire_R_0; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_10;
  reg  output_fire_R_1; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_11;
  reg  output_fire_R_2; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_12;
  reg  output_fire_R_3; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_13;
  reg  output_fire_R_4; // @[BasicBlock.scala 227:48]
  reg [31:0] _RAND_14;
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[BasicBlock.scala 232:36]
  wire [4:0] in_task_ID; // @[BasicBlock.scala 239:34]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[BasicBlock.scala 244:28]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BasicBlock.scala 244:28]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[BasicBlock.scala 244:28]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_10; // @[BasicBlock.scala 244:28]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_12; // @[BasicBlock.scala 244:28]
  wire  out_fire_mask_0; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_1; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_2; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_3; // @[BasicBlock.scala 256:85]
  wire  out_fire_mask_4; // @[BasicBlock.scala 256:85]
  reg  state; // @[BasicBlock.scala 292:22]
  reg [31:0] _RAND_15;
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_33; // @[BasicBlock.scala 309:81]
  wire  _T_34; // @[BasicBlock.scala 309:81]
  wire  _T_35; // @[BasicBlock.scala 309:81]
  wire  _T_36; // @[BasicBlock.scala 309:81]
  wire  _T_37; // @[BasicBlock.scala 309:81]
  wire  _T_38; // @[BasicBlock.scala 315:19]
  wire  _T_39; // @[BasicBlock.scala 315:19]
  wire  _GEN_14; // @[BasicBlock.scala 304:8]
  wire  _GEN_15; // @[BasicBlock.scala 304:8]
  wire  _GEN_16; // @[BasicBlock.scala 304:8]
  wire  _GEN_17; // @[BasicBlock.scala 304:8]
  wire  _GEN_18; // @[BasicBlock.scala 304:8]
  wire  _GEN_24; // @[BasicBlock.scala 304:8]
  wire  _T_43; // @[BasicBlock.scala 328:35]
  wire  _T_44; // @[BasicBlock.scala 328:35]
  wire  _T_45; // @[BasicBlock.scala 328:35]
  wire  _T_46; // @[BasicBlock.scala 328:35]
  wire  _GEN_62; // @[BasicBlock.scala 315:19]
  wire  _GEN_63; // @[BasicBlock.scala 315:19]
  wire  _GEN_65; // @[BasicBlock.scala 320:19]
  wire  _GEN_66; // @[BasicBlock.scala 320:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_7 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_7 | in_data_valid_R_0; // @[BasicBlock.scala 232:36]
  assign in_task_ID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 239:34]
  assign _T_8 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_8 | output_fire_R_0; // @[BasicBlock.scala 244:28]
  assign _T_9 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_9 | output_fire_R_1; // @[BasicBlock.scala 244:28]
  assign _T_10 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 | output_fire_R_2; // @[BasicBlock.scala 244:28]
  assign _T_11 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_10 = _T_11 | output_fire_R_3; // @[BasicBlock.scala 244:28]
  assign _T_12 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_12 = _T_12 | output_fire_R_4; // @[BasicBlock.scala 244:28]
  assign out_fire_mask_0 = output_fire_R_0 | _T_8; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_1 = output_fire_R_1 | _T_9; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_2 = output_fire_R_2 | _T_10; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_3 = output_fire_R_3 | _T_11; // @[BasicBlock.scala 256:85]
  assign out_fire_mask_4 = output_fire_R_4 | _T_12; // @[BasicBlock.scala 256:85]
  assign _T_27 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_33 = _T_8 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_34 = _T_9 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_35 = _T_10 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_36 = _T_11 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_37 = _T_12 ^ 1'h1; // @[BasicBlock.scala 309:81]
  assign _T_38 = $unsigned(reset); // @[BasicBlock.scala 315:19]
  assign _T_39 = _T_38 == 1'h0; // @[BasicBlock.scala 315:19]
  assign _GEN_14 = _GEN_3 | output_valid_R_0; // @[BasicBlock.scala 304:8]
  assign _GEN_15 = _GEN_3 | output_valid_R_1; // @[BasicBlock.scala 304:8]
  assign _GEN_16 = _GEN_3 | output_valid_R_2; // @[BasicBlock.scala 304:8]
  assign _GEN_17 = _GEN_3 | output_valid_R_3; // @[BasicBlock.scala 304:8]
  assign _GEN_18 = _GEN_3 | output_valid_R_4; // @[BasicBlock.scala 304:8]
  assign _GEN_24 = _GEN_3 | state; // @[BasicBlock.scala 304:8]
  assign _T_43 = out_fire_mask_0 & out_fire_mask_1; // @[BasicBlock.scala 328:35]
  assign _T_44 = _T_43 & out_fire_mask_2; // @[BasicBlock.scala 328:35]
  assign _T_45 = _T_44 & out_fire_mask_3; // @[BasicBlock.scala 328:35]
  assign _T_46 = _T_45 & out_fire_mask_4; // @[BasicBlock.scala 328:35]
  assign io_predicateIn_0_ready = ~ in_data_valid_R_0; // @[BasicBlock.scala 231:29]
  assign io_Out_0_valid = _T_27 ? _GEN_14 : output_valid_R_0; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_0_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_1_valid = _T_27 ? _GEN_15 : output_valid_R_1; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_1_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_2_valid = _T_27 ? _GEN_16 : output_valid_R_2; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_2_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_2_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_3_valid = _T_27 ? _GEN_17 : output_valid_R_3; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_3_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_3_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign io_Out_4_valid = _T_27 ? _GEN_18 : output_valid_R_4; // @[BasicBlock.scala 287:21 BasicBlock.scala 306:34]
  assign io_Out_4_bits_taskID = io_predicateIn_0_bits_taskID | in_data_R_0_taskID; // @[BasicBlock.scala 282:22]
  assign io_Out_4_bits_control = _T_7 ? io_predicateIn_0_bits_control : in_data_R_0_control; // @[BasicBlock.scala 282:22]
  assign _GEN_62 = _T_27 & _GEN_3; // @[BasicBlock.scala 315:19]
  assign _GEN_63 = _GEN_62 & in_data_R_0_control; // @[BasicBlock.scala 315:19]
  assign _GEN_65 = in_data_R_0_control == 1'h0; // @[BasicBlock.scala 320:19]
  assign _GEN_66 = _GEN_62 & _GEN_65; // @[BasicBlock.scala 320:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_0_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_R_0_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  output_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_valid_R_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_valid_R_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  output_valid_R_4 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_fire_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_fire_R_1 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_fire_R_2 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  output_fire_R_3 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  output_fire_R_4 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  state = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_0_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_7) begin
          in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_46) begin
            in_data_R_0_taskID <= 5'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_taskID <= io_predicateIn_0_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      in_data_R_0_control <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_7) begin
          in_data_R_0_control <= io_predicateIn_0_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_46) begin
            in_data_R_0_control <= 1'h0;
          end else begin
            if (_T_7) begin
              in_data_R_0_control <= io_predicateIn_0_bits_control;
            end
          end
        end else begin
          if (_T_7) begin
            in_data_R_0_control <= io_predicateIn_0_bits_control;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_27) begin
        in_data_valid_R_0 <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_46) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_3;
          end
        end else begin
          in_data_valid_R_0 <= _GEN_3;
        end
      end
    end
    if (reset) begin
      output_R_taskID <= 5'h0;
    end else begin
      output_R_taskID <= in_task_ID;
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_0 <= _T_33;
        end else begin
          if (_T_8) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          output_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_1 <= _T_34;
        end else begin
          if (_T_9) begin
            output_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_9) begin
          output_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_2 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_2 <= _T_35;
        end else begin
          if (_T_10) begin
            output_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_10) begin
          output_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_3 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_3 <= _T_36;
        end else begin
          if (_T_11) begin
            output_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_11) begin
          output_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_valid_R_4 <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_GEN_3) begin
          output_valid_R_4 <= _T_37;
        end else begin
          if (_T_12) begin
            output_valid_R_4 <= 1'h0;
          end
        end
      end else begin
        if (_T_12) begin
          output_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      output_fire_R_0 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_0 <= _GEN_4;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_0 <= 1'h0;
          end else begin
            output_fire_R_0 <= _GEN_4;
          end
        end else begin
          output_fire_R_0 <= _GEN_4;
        end
      end
    end
    if (reset) begin
      output_fire_R_1 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_1 <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_1 <= 1'h0;
          end else begin
            output_fire_R_1 <= _GEN_6;
          end
        end else begin
          output_fire_R_1 <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_fire_R_2 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_2 <= _GEN_8;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_2 <= 1'h0;
          end else begin
            output_fire_R_2 <= _GEN_8;
          end
        end else begin
          output_fire_R_2 <= _GEN_8;
        end
      end
    end
    if (reset) begin
      output_fire_R_3 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_3 <= _GEN_10;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_3 <= 1'h0;
          end else begin
            output_fire_R_3 <= _GEN_10;
          end
        end else begin
          output_fire_R_3 <= _GEN_10;
        end
      end
    end
    if (reset) begin
      output_fire_R_4 <= 1'h0;
    end else begin
      if (_T_27) begin
        output_fire_R_4 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_46) begin
            output_fire_R_4 <= 1'h0;
          end else begin
            output_fire_R_4 <= _GEN_12;
          end
        end else begin
          output_fire_R_4 <= _GEN_12;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_27) begin
        state <= _GEN_24;
      end else begin
        if (state) begin
          if (_T_46) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [BB]   bb_for_cond_cleanup113: Output [T] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 315:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_66 & _T_39) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [BB]   bb_for_cond_cleanup113: Output [F] fired @ %d\n",output_R_taskID,value); // @[BasicBlock.scala 320:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BasicBlockNode_1(
  input        clock,
  input        reset,
  input        io_MaskBB_0_ready,
  output       io_MaskBB_0_valid,
  output [1:0] io_MaskBB_0_bits,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  input        io_Out_1_ready,
  output       io_Out_1_valid,
  output [4:0] io_Out_1_bits_taskID,
  input        io_Out_2_ready,
  output       io_Out_2_valid,
  output [4:0] io_Out_2_bits_taskID,
  input        io_Out_3_ready,
  output       io_Out_3_valid,
  output [4:0] io_Out_3_bits_taskID,
  input        io_Out_4_ready,
  output       io_Out_4_valid,
  output [4:0] io_Out_4_bits_taskID,
  input        io_Out_5_ready,
  output       io_Out_5_valid,
  output [4:0] io_Out_5_bits_taskID,
  input        io_Out_6_ready,
  output       io_Out_6_valid,
  output [4:0] io_Out_6_bits_taskID,
  input        io_Out_7_ready,
  output       io_Out_7_valid,
  output [4:0] io_Out_7_bits_taskID,
  input        io_Out_8_ready,
  output       io_Out_8_valid,
  output [4:0] io_Out_8_bits_taskID,
  input        io_Out_9_ready,
  output       io_Out_9_valid,
  output [4:0] io_Out_9_bits_taskID,
  input        io_Out_10_ready,
  output       io_Out_10_valid,
  output [4:0] io_Out_10_bits_taskID,
  input        io_Out_11_ready,
  output       io_Out_11_valid,
  output       io_Out_11_bits_control,
  input        io_Out_12_ready,
  output       io_Out_12_valid,
  output [4:0] io_Out_12_bits_taskID,
  output       io_Out_12_bits_control,
  input        io_Out_13_ready,
  output       io_Out_13_valid,
  output [4:0] io_Out_13_bits_taskID,
  output       io_Out_13_bits_control,
  input        io_Out_14_ready,
  output       io_Out_14_valid,
  output [4:0] io_Out_14_bits_taskID,
  output       io_Out_14_bits_control,
  input        io_Out_15_ready,
  output       io_Out_15_valid,
  output [4:0] io_Out_15_bits_taskID,
  output       io_Out_15_bits_control,
  input        io_Out_16_ready,
  output       io_Out_16_valid,
  output [4:0] io_Out_16_bits_taskID,
  output       io_Out_16_bits_control,
  input        io_Out_17_ready,
  output       io_Out_17_valid,
  output [4:0] io_Out_17_bits_taskID,
  output       io_Out_17_bits_control,
  input        io_Out_18_ready,
  output       io_Out_18_valid,
  output [4:0] io_Out_18_bits_taskID,
  output       io_Out_18_bits_control,
  input        io_Out_19_ready,
  output       io_Out_19_valid,
  output [4:0] io_Out_19_bits_taskID,
  output       io_Out_19_bits_control,
  input        io_Out_20_ready,
  output       io_Out_20_valid,
  output [4:0] io_Out_20_bits_taskID,
  output       io_Out_20_bits_control,
  input        io_Out_21_ready,
  output       io_Out_21_valid,
  output [4:0] io_Out_21_bits_taskID,
  input        io_Out_22_ready,
  output       io_Out_22_valid,
  output [4:0] io_Out_22_bits_taskID,
  output       io_Out_22_bits_control,
  input        io_Out_23_ready,
  output       io_Out_23_valid,
  output [4:0] io_Out_23_bits_taskID,
  output       io_Out_23_bits_control,
  input        io_Out_24_ready,
  output       io_Out_24_valid,
  output [4:0] io_Out_24_bits_taskID,
  output       io_Out_24_bits_control,
  input        io_Out_25_ready,
  output       io_Out_25_valid,
  output [4:0] io_Out_25_bits_taskID,
  output       io_Out_25_bits_control,
  input        io_Out_26_ready,
  output       io_Out_26_valid,
  output [4:0] io_Out_26_bits_taskID,
  output       io_Out_26_bits_control,
  input        io_Out_27_ready,
  output       io_Out_27_valid,
  output [4:0] io_Out_27_bits_taskID,
  output       io_Out_27_bits_control,
  input        io_Out_28_ready,
  output       io_Out_28_valid,
  output [4:0] io_Out_28_bits_taskID,
  output       io_Out_28_bits_control,
  input        io_Out_29_ready,
  output       io_Out_29_valid,
  output [4:0] io_Out_29_bits_taskID,
  input        io_Out_30_ready,
  output       io_Out_30_valid,
  output [4:0] io_Out_30_bits_taskID,
  output       io_Out_30_bits_control,
  input        io_Out_31_ready,
  output       io_Out_31_valid,
  output [4:0] io_Out_31_bits_taskID,
  output       io_Out_31_bits_control,
  input        io_Out_32_ready,
  output       io_Out_32_valid,
  output [4:0] io_Out_32_bits_taskID,
  output       io_Out_32_bits_control,
  input        io_Out_33_ready,
  output       io_Out_33_valid,
  output [4:0] io_Out_33_bits_taskID,
  output       io_Out_33_bits_control,
  input        io_Out_34_ready,
  output       io_Out_34_valid,
  output [4:0] io_Out_34_bits_taskID,
  output       io_Out_34_bits_control,
  input        io_Out_35_ready,
  output       io_Out_35_valid,
  output [4:0] io_Out_35_bits_taskID,
  output       io_Out_35_bits_control,
  input        io_Out_36_ready,
  output       io_Out_36_valid,
  output [4:0] io_Out_36_bits_taskID,
  output       io_Out_36_bits_control,
  input        io_Out_37_ready,
  output       io_Out_37_valid,
  output [4:0] io_Out_37_bits_taskID,
  input        io_Out_38_ready,
  output       io_Out_38_valid,
  output [4:0] io_Out_38_bits_taskID,
  output       io_Out_38_bits_control,
  input        io_Out_39_ready,
  output       io_Out_39_valid,
  output [4:0] io_Out_39_bits_taskID,
  output       io_Out_39_bits_control,
  input        io_Out_40_ready,
  output       io_Out_40_valid,
  output [4:0] io_Out_40_bits_taskID,
  output       io_Out_40_bits_control,
  input        io_Out_41_ready,
  output       io_Out_41_valid,
  output [4:0] io_Out_41_bits_taskID,
  output       io_Out_41_bits_control,
  input        io_Out_42_ready,
  output       io_Out_42_valid,
  output [4:0] io_Out_42_bits_taskID,
  output       io_Out_42_bits_control,
  input        io_Out_43_ready,
  output       io_Out_43_valid,
  output [4:0] io_Out_43_bits_taskID,
  output       io_Out_43_bits_control,
  input        io_Out_44_ready,
  output       io_Out_44_valid,
  output [4:0] io_Out_44_bits_taskID,
  output       io_Out_44_bits_control,
  input        io_Out_45_ready,
  output       io_Out_45_valid,
  output [4:0] io_Out_45_bits_taskID,
  output       io_Out_45_bits_control,
  input        io_Out_46_ready,
  output       io_Out_46_valid,
  output [4:0] io_Out_46_bits_taskID,
  input        io_Out_47_ready,
  output       io_Out_47_valid,
  output [4:0] io_Out_47_bits_taskID,
  output       io_Out_47_bits_control,
  input        io_Out_48_ready,
  output       io_Out_48_valid,
  output [4:0] io_Out_48_bits_taskID,
  output       io_Out_48_bits_control,
  input        io_Out_49_ready,
  output       io_Out_49_valid,
  output [4:0] io_Out_49_bits_taskID,
  output       io_Out_49_bits_control,
  input        io_Out_50_ready,
  output       io_Out_50_valid,
  output [4:0] io_Out_50_bits_taskID,
  output       io_Out_50_bits_control,
  input        io_Out_51_ready,
  output       io_Out_51_valid,
  output [4:0] io_Out_51_bits_taskID,
  output       io_Out_51_bits_control,
  input        io_Out_52_ready,
  output       io_Out_52_valid,
  output [4:0] io_Out_52_bits_taskID,
  output       io_Out_52_bits_control,
  input        io_Out_53_ready,
  output       io_Out_53_valid,
  output [4:0] io_Out_53_bits_taskID,
  output       io_Out_53_bits_control,
  input        io_Out_54_ready,
  output       io_Out_54_valid,
  output [4:0] io_Out_54_bits_taskID,
  input        io_Out_55_ready,
  output       io_Out_55_valid,
  output [4:0] io_Out_55_bits_taskID,
  output       io_Out_55_bits_control,
  input        io_Out_56_ready,
  output       io_Out_56_valid,
  output [4:0] io_Out_56_bits_taskID,
  output       io_Out_56_bits_control,
  input        io_Out_57_ready,
  output       io_Out_57_valid,
  output [4:0] io_Out_57_bits_taskID,
  output       io_Out_57_bits_control,
  input        io_Out_58_ready,
  output       io_Out_58_valid,
  output [4:0] io_Out_58_bits_taskID,
  output       io_Out_58_bits_control,
  input        io_Out_59_ready,
  output       io_Out_59_valid,
  output [4:0] io_Out_59_bits_taskID,
  output       io_Out_59_bits_control,
  input        io_Out_60_ready,
  output       io_Out_60_valid,
  output [4:0] io_Out_60_bits_taskID,
  output       io_Out_60_bits_control,
  input        io_Out_61_ready,
  output       io_Out_61_valid,
  output [4:0] io_Out_61_bits_taskID,
  output       io_Out_61_bits_control,
  input        io_Out_62_ready,
  output       io_Out_62_valid,
  output [4:0] io_Out_62_bits_taskID,
  input        io_Out_63_ready,
  output       io_Out_63_valid,
  output [4:0] io_Out_63_bits_taskID,
  output       io_Out_63_bits_control,
  input        io_Out_64_ready,
  output       io_Out_64_valid,
  output [4:0] io_Out_64_bits_taskID,
  output       io_Out_64_bits_control,
  input        io_Out_65_ready,
  output       io_Out_65_valid,
  output [4:0] io_Out_65_bits_taskID,
  output       io_Out_65_bits_control,
  input        io_Out_66_ready,
  output       io_Out_66_valid,
  output [4:0] io_Out_66_bits_taskID,
  output       io_Out_66_bits_control,
  input        io_Out_67_ready,
  output       io_Out_67_valid,
  output [4:0] io_Out_67_bits_taskID,
  output       io_Out_67_bits_control,
  input        io_Out_68_ready,
  output       io_Out_68_valid,
  output [4:0] io_Out_68_bits_taskID,
  output       io_Out_68_bits_control,
  input        io_Out_69_ready,
  output       io_Out_69_valid,
  output [4:0] io_Out_69_bits_taskID,
  output       io_Out_69_bits_control,
  input        io_Out_70_ready,
  output       io_Out_70_valid,
  output [4:0] io_Out_70_bits_taskID,
  input        io_Out_71_ready,
  output       io_Out_71_valid,
  output [4:0] io_Out_71_bits_taskID,
  output       io_Out_71_bits_control,
  input        io_Out_72_ready,
  output       io_Out_72_valid,
  output [4:0] io_Out_72_bits_taskID,
  output       io_Out_72_bits_control,
  input        io_Out_73_ready,
  output       io_Out_73_valid,
  output [4:0] io_Out_73_bits_taskID,
  output       io_Out_73_bits_control,
  input        io_Out_74_ready,
  output       io_Out_74_valid,
  output [4:0] io_Out_74_bits_taskID,
  output       io_Out_74_bits_control,
  input        io_Out_75_ready,
  output       io_Out_75_valid,
  output [4:0] io_Out_75_bits_taskID,
  output       io_Out_75_bits_control,
  input        io_Out_76_ready,
  output       io_Out_76_valid,
  output [4:0] io_Out_76_bits_taskID,
  output       io_Out_76_bits_control,
  input        io_Out_77_ready,
  output       io_Out_77_valid,
  output [4:0] io_Out_77_bits_taskID,
  output       io_Out_77_bits_control,
  input        io_Out_78_ready,
  output       io_Out_78_valid,
  output [4:0] io_Out_78_bits_taskID,
  input        io_Out_79_ready,
  output       io_Out_79_valid,
  output [4:0] io_Out_79_bits_taskID,
  output       io_Out_79_bits_control,
  input        io_Out_80_ready,
  output       io_Out_80_valid,
  output [4:0] io_Out_80_bits_taskID,
  output       io_Out_80_bits_control,
  input        io_Out_81_ready,
  output       io_Out_81_valid,
  output [4:0] io_Out_81_bits_taskID,
  output       io_Out_81_bits_control,
  input        io_Out_82_ready,
  output       io_Out_82_valid,
  output [4:0] io_Out_82_bits_taskID,
  output       io_Out_82_bits_control,
  input        io_Out_83_ready,
  output       io_Out_83_valid,
  output [4:0] io_Out_83_bits_taskID,
  output       io_Out_83_bits_control,
  input        io_Out_84_ready,
  output       io_Out_84_valid,
  output [4:0] io_Out_84_bits_taskID,
  output       io_Out_84_bits_control,
  input        io_Out_85_ready,
  output       io_Out_85_valid,
  output [4:0] io_Out_85_bits_taskID,
  output       io_Out_85_bits_control,
  input        io_Out_86_ready,
  output       io_Out_86_valid,
  output [4:0] io_Out_86_bits_taskID,
  input        io_Out_87_ready,
  output       io_Out_87_valid,
  output [4:0] io_Out_87_bits_taskID,
  output       io_Out_87_bits_control,
  input        io_Out_88_ready,
  output       io_Out_88_valid,
  output [4:0] io_Out_88_bits_taskID,
  output       io_Out_88_bits_control,
  input        io_Out_89_ready,
  output       io_Out_89_valid,
  output [4:0] io_Out_89_bits_taskID,
  output       io_Out_89_bits_control,
  input        io_Out_90_ready,
  output       io_Out_90_valid,
  output [4:0] io_Out_90_bits_taskID,
  output       io_Out_90_bits_control,
  input        io_Out_91_ready,
  output       io_Out_91_valid,
  output [4:0] io_Out_91_bits_taskID,
  output       io_Out_91_bits_control,
  input        io_Out_92_ready,
  output       io_Out_92_valid,
  output [4:0] io_Out_92_bits_taskID,
  output       io_Out_92_bits_control,
  output       io_predicateIn_0_ready,
  input        io_predicateIn_0_valid,
  input  [4:0] io_predicateIn_0_bits_taskID,
  input        io_predicateIn_0_bits_control,
  output       io_predicateIn_1_ready,
  input        io_predicateIn_1_valid,
  input  [4:0] io_predicateIn_1_bits_taskID,
  input        io_predicateIn_1_bits_control
);
  reg  out_ready_R_0; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_0;
  reg  out_ready_R_1; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_1;
  reg  out_ready_R_2; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_2;
  reg  out_ready_R_3; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_3;
  reg  out_ready_R_4; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_4;
  reg  out_ready_R_5; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_5;
  reg  out_ready_R_6; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_6;
  reg  out_ready_R_7; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_7;
  reg  out_ready_R_8; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_8;
  reg  out_ready_R_9; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_9;
  reg  out_ready_R_10; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_10;
  reg  out_ready_R_11; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_11;
  reg  out_ready_R_12; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_12;
  reg  out_ready_R_13; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_13;
  reg  out_ready_R_14; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_14;
  reg  out_ready_R_15; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_15;
  reg  out_ready_R_16; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_16;
  reg  out_ready_R_17; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_17;
  reg  out_ready_R_18; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_18;
  reg  out_ready_R_19; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_19;
  reg  out_ready_R_20; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_20;
  reg  out_ready_R_21; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_21;
  reg  out_ready_R_22; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_22;
  reg  out_ready_R_23; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_23;
  reg  out_ready_R_24; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_24;
  reg  out_ready_R_25; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_25;
  reg  out_ready_R_26; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_26;
  reg  out_ready_R_27; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_27;
  reg  out_ready_R_28; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_28;
  reg  out_ready_R_29; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_29;
  reg  out_ready_R_30; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_30;
  reg  out_ready_R_31; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_31;
  reg  out_ready_R_32; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_32;
  reg  out_ready_R_33; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_33;
  reg  out_ready_R_34; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_34;
  reg  out_ready_R_35; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_35;
  reg  out_ready_R_36; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_36;
  reg  out_ready_R_37; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_37;
  reg  out_ready_R_38; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_38;
  reg  out_ready_R_39; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_39;
  reg  out_ready_R_40; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_40;
  reg  out_ready_R_41; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_41;
  reg  out_ready_R_42; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_42;
  reg  out_ready_R_43; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_43;
  reg  out_ready_R_44; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_44;
  reg  out_ready_R_45; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_45;
  reg  out_ready_R_46; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_46;
  reg  out_ready_R_47; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_47;
  reg  out_ready_R_48; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_48;
  reg  out_ready_R_49; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_49;
  reg  out_ready_R_50; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_50;
  reg  out_ready_R_51; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_51;
  reg  out_ready_R_52; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_52;
  reg  out_ready_R_53; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_53;
  reg  out_ready_R_54; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_54;
  reg  out_ready_R_55; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_55;
  reg  out_ready_R_56; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_56;
  reg  out_ready_R_57; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_57;
  reg  out_ready_R_58; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_58;
  reg  out_ready_R_59; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_59;
  reg  out_ready_R_60; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_60;
  reg  out_ready_R_61; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_61;
  reg  out_ready_R_62; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_62;
  reg  out_ready_R_63; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_63;
  reg  out_ready_R_64; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_64;
  reg  out_ready_R_65; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_65;
  reg  out_ready_R_66; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_66;
  reg  out_ready_R_67; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_67;
  reg  out_ready_R_68; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_68;
  reg  out_ready_R_69; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_69;
  reg  out_ready_R_70; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_70;
  reg  out_ready_R_71; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_71;
  reg  out_ready_R_72; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_72;
  reg  out_ready_R_73; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_73;
  reg  out_ready_R_74; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_74;
  reg  out_ready_R_75; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_75;
  reg  out_ready_R_76; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_76;
  reg  out_ready_R_77; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_77;
  reg  out_ready_R_78; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_78;
  reg  out_ready_R_79; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_79;
  reg  out_ready_R_80; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_80;
  reg  out_ready_R_81; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_81;
  reg  out_ready_R_82; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_82;
  reg  out_ready_R_83; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_83;
  reg  out_ready_R_84; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_84;
  reg  out_ready_R_85; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_85;
  reg  out_ready_R_86; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_86;
  reg  out_ready_R_87; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_87;
  reg  out_ready_R_88; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_88;
  reg  out_ready_R_89; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_89;
  reg  out_ready_R_90; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_90;
  reg  out_ready_R_91; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_91;
  reg  out_ready_R_92; // @[HandShaking.scala 702:28]
  reg [31:0] _RAND_92;
  reg  out_valid_R_0; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_93;
  reg  out_valid_R_1; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_94;
  reg  out_valid_R_2; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_95;
  reg  out_valid_R_3; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_96;
  reg  out_valid_R_4; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_97;
  reg  out_valid_R_5; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_98;
  reg  out_valid_R_6; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_99;
  reg  out_valid_R_7; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_100;
  reg  out_valid_R_8; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_101;
  reg  out_valid_R_9; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_102;
  reg  out_valid_R_10; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_103;
  reg  out_valid_R_11; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_104;
  reg  out_valid_R_12; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_105;
  reg  out_valid_R_13; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_106;
  reg  out_valid_R_14; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_107;
  reg  out_valid_R_15; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_108;
  reg  out_valid_R_16; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_109;
  reg  out_valid_R_17; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_110;
  reg  out_valid_R_18; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_111;
  reg  out_valid_R_19; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_112;
  reg  out_valid_R_20; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_113;
  reg  out_valid_R_21; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_114;
  reg  out_valid_R_22; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_115;
  reg  out_valid_R_23; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_116;
  reg  out_valid_R_24; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_117;
  reg  out_valid_R_25; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_118;
  reg  out_valid_R_26; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_119;
  reg  out_valid_R_27; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_120;
  reg  out_valid_R_28; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_121;
  reg  out_valid_R_29; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_122;
  reg  out_valid_R_30; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_123;
  reg  out_valid_R_31; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_124;
  reg  out_valid_R_32; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_125;
  reg  out_valid_R_33; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_126;
  reg  out_valid_R_34; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_127;
  reg  out_valid_R_35; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_128;
  reg  out_valid_R_36; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_129;
  reg  out_valid_R_37; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_130;
  reg  out_valid_R_38; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_131;
  reg  out_valid_R_39; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_132;
  reg  out_valid_R_40; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_133;
  reg  out_valid_R_41; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_134;
  reg  out_valid_R_42; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_135;
  reg  out_valid_R_43; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_136;
  reg  out_valid_R_44; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_137;
  reg  out_valid_R_45; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_138;
  reg  out_valid_R_46; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_139;
  reg  out_valid_R_47; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_140;
  reg  out_valid_R_48; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_141;
  reg  out_valid_R_49; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_142;
  reg  out_valid_R_50; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_143;
  reg  out_valid_R_51; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_144;
  reg  out_valid_R_52; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_145;
  reg  out_valid_R_53; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_146;
  reg  out_valid_R_54; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_147;
  reg  out_valid_R_55; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_148;
  reg  out_valid_R_56; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_149;
  reg  out_valid_R_57; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_150;
  reg  out_valid_R_58; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_151;
  reg  out_valid_R_59; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_152;
  reg  out_valid_R_60; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_153;
  reg  out_valid_R_61; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_154;
  reg  out_valid_R_62; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_155;
  reg  out_valid_R_63; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_156;
  reg  out_valid_R_64; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_157;
  reg  out_valid_R_65; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_158;
  reg  out_valid_R_66; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_159;
  reg  out_valid_R_67; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_160;
  reg  out_valid_R_68; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_161;
  reg  out_valid_R_69; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_162;
  reg  out_valid_R_70; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_163;
  reg  out_valid_R_71; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_164;
  reg  out_valid_R_72; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_165;
  reg  out_valid_R_73; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_166;
  reg  out_valid_R_74; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_167;
  reg  out_valid_R_75; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_168;
  reg  out_valid_R_76; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_169;
  reg  out_valid_R_77; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_170;
  reg  out_valid_R_78; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_171;
  reg  out_valid_R_79; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_172;
  reg  out_valid_R_80; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_173;
  reg  out_valid_R_81; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_174;
  reg  out_valid_R_82; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_175;
  reg  out_valid_R_83; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_176;
  reg  out_valid_R_84; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_177;
  reg  out_valid_R_85; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_178;
  reg  out_valid_R_86; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_179;
  reg  out_valid_R_87; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_180;
  reg  out_valid_R_88; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_181;
  reg  out_valid_R_89; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_182;
  reg  out_valid_R_90; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_183;
  reg  out_valid_R_91; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_184;
  reg  out_valid_R_92; // @[HandShaking.scala 703:28]
  reg [31:0] _RAND_185;
  reg  mask_valid_R_0; // @[HandShaking.scala 707:46]
  reg [31:0] _RAND_186;
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _GEN_1; // @[HandShaking.scala 716:29]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _GEN_3; // @[HandShaking.scala 716:29]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[HandShaking.scala 716:29]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[HandShaking.scala 716:29]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[HandShaking.scala 716:29]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[HandShaking.scala 716:29]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[HandShaking.scala 716:29]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[HandShaking.scala 716:29]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[HandShaking.scala 716:29]
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[HandShaking.scala 716:29]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_21; // @[HandShaking.scala 716:29]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_23; // @[HandShaking.scala 716:29]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_25; // @[HandShaking.scala 716:29]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_27; // @[HandShaking.scala 716:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_29; // @[HandShaking.scala 716:29]
  wire  _T_17; // @[Decoupled.scala 40:37]
  wire  _GEN_31; // @[HandShaking.scala 716:29]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_33; // @[HandShaking.scala 716:29]
  wire  _T_19; // @[Decoupled.scala 40:37]
  wire  _GEN_35; // @[HandShaking.scala 716:29]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_37; // @[HandShaking.scala 716:29]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_39; // @[HandShaking.scala 716:29]
  wire  _T_22; // @[Decoupled.scala 40:37]
  wire  _GEN_41; // @[HandShaking.scala 716:29]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _GEN_43; // @[HandShaking.scala 716:29]
  wire  _T_24; // @[Decoupled.scala 40:37]
  wire  _GEN_45; // @[HandShaking.scala 716:29]
  wire  _T_25; // @[Decoupled.scala 40:37]
  wire  _GEN_47; // @[HandShaking.scala 716:29]
  wire  _T_26; // @[Decoupled.scala 40:37]
  wire  _GEN_49; // @[HandShaking.scala 716:29]
  wire  _T_27; // @[Decoupled.scala 40:37]
  wire  _GEN_51; // @[HandShaking.scala 716:29]
  wire  _T_28; // @[Decoupled.scala 40:37]
  wire  _GEN_53; // @[HandShaking.scala 716:29]
  wire  _T_29; // @[Decoupled.scala 40:37]
  wire  _GEN_55; // @[HandShaking.scala 716:29]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_57; // @[HandShaking.scala 716:29]
  wire  _T_31; // @[Decoupled.scala 40:37]
  wire  _GEN_59; // @[HandShaking.scala 716:29]
  wire  _T_32; // @[Decoupled.scala 40:37]
  wire  _GEN_61; // @[HandShaking.scala 716:29]
  wire  _T_33; // @[Decoupled.scala 40:37]
  wire  _GEN_63; // @[HandShaking.scala 716:29]
  wire  _T_34; // @[Decoupled.scala 40:37]
  wire  _GEN_65; // @[HandShaking.scala 716:29]
  wire  _T_35; // @[Decoupled.scala 40:37]
  wire  _GEN_67; // @[HandShaking.scala 716:29]
  wire  _T_36; // @[Decoupled.scala 40:37]
  wire  _GEN_69; // @[HandShaking.scala 716:29]
  wire  _T_37; // @[Decoupled.scala 40:37]
  wire  _GEN_71; // @[HandShaking.scala 716:29]
  wire  _T_38; // @[Decoupled.scala 40:37]
  wire  _GEN_73; // @[HandShaking.scala 716:29]
  wire  _T_39; // @[Decoupled.scala 40:37]
  wire  _GEN_75; // @[HandShaking.scala 716:29]
  wire  _T_40; // @[Decoupled.scala 40:37]
  wire  _GEN_77; // @[HandShaking.scala 716:29]
  wire  _T_41; // @[Decoupled.scala 40:37]
  wire  _GEN_79; // @[HandShaking.scala 716:29]
  wire  _T_42; // @[Decoupled.scala 40:37]
  wire  _GEN_81; // @[HandShaking.scala 716:29]
  wire  _T_43; // @[Decoupled.scala 40:37]
  wire  _GEN_83; // @[HandShaking.scala 716:29]
  wire  _T_44; // @[Decoupled.scala 40:37]
  wire  _GEN_85; // @[HandShaking.scala 716:29]
  wire  _T_45; // @[Decoupled.scala 40:37]
  wire  _GEN_87; // @[HandShaking.scala 716:29]
  wire  _T_46; // @[Decoupled.scala 40:37]
  wire  _GEN_89; // @[HandShaking.scala 716:29]
  wire  _T_47; // @[Decoupled.scala 40:37]
  wire  _GEN_91; // @[HandShaking.scala 716:29]
  wire  _T_48; // @[Decoupled.scala 40:37]
  wire  _GEN_93; // @[HandShaking.scala 716:29]
  wire  _T_49; // @[Decoupled.scala 40:37]
  wire  _GEN_95; // @[HandShaking.scala 716:29]
  wire  _T_50; // @[Decoupled.scala 40:37]
  wire  _GEN_97; // @[HandShaking.scala 716:29]
  wire  _T_51; // @[Decoupled.scala 40:37]
  wire  _GEN_99; // @[HandShaking.scala 716:29]
  wire  _T_52; // @[Decoupled.scala 40:37]
  wire  _GEN_101; // @[HandShaking.scala 716:29]
  wire  _T_53; // @[Decoupled.scala 40:37]
  wire  _GEN_103; // @[HandShaking.scala 716:29]
  wire  _T_54; // @[Decoupled.scala 40:37]
  wire  _GEN_105; // @[HandShaking.scala 716:29]
  wire  _T_55; // @[Decoupled.scala 40:37]
  wire  _GEN_107; // @[HandShaking.scala 716:29]
  wire  _T_56; // @[Decoupled.scala 40:37]
  wire  _GEN_109; // @[HandShaking.scala 716:29]
  wire  _T_57; // @[Decoupled.scala 40:37]
  wire  _GEN_111; // @[HandShaking.scala 716:29]
  wire  _T_58; // @[Decoupled.scala 40:37]
  wire  _GEN_113; // @[HandShaking.scala 716:29]
  wire  _T_59; // @[Decoupled.scala 40:37]
  wire  _GEN_115; // @[HandShaking.scala 716:29]
  wire  _T_60; // @[Decoupled.scala 40:37]
  wire  _GEN_117; // @[HandShaking.scala 716:29]
  wire  _T_61; // @[Decoupled.scala 40:37]
  wire  _GEN_119; // @[HandShaking.scala 716:29]
  wire  _T_62; // @[Decoupled.scala 40:37]
  wire  _GEN_121; // @[HandShaking.scala 716:29]
  wire  _T_63; // @[Decoupled.scala 40:37]
  wire  _GEN_123; // @[HandShaking.scala 716:29]
  wire  _T_64; // @[Decoupled.scala 40:37]
  wire  _GEN_125; // @[HandShaking.scala 716:29]
  wire  _T_65; // @[Decoupled.scala 40:37]
  wire  _GEN_127; // @[HandShaking.scala 716:29]
  wire  _T_66; // @[Decoupled.scala 40:37]
  wire  _GEN_129; // @[HandShaking.scala 716:29]
  wire  _T_67; // @[Decoupled.scala 40:37]
  wire  _GEN_131; // @[HandShaking.scala 716:29]
  wire  _T_68; // @[Decoupled.scala 40:37]
  wire  _GEN_133; // @[HandShaking.scala 716:29]
  wire  _T_69; // @[Decoupled.scala 40:37]
  wire  _GEN_135; // @[HandShaking.scala 716:29]
  wire  _T_70; // @[Decoupled.scala 40:37]
  wire  _GEN_137; // @[HandShaking.scala 716:29]
  wire  _T_71; // @[Decoupled.scala 40:37]
  wire  _GEN_139; // @[HandShaking.scala 716:29]
  wire  _T_72; // @[Decoupled.scala 40:37]
  wire  _GEN_141; // @[HandShaking.scala 716:29]
  wire  _T_73; // @[Decoupled.scala 40:37]
  wire  _GEN_143; // @[HandShaking.scala 716:29]
  wire  _T_74; // @[Decoupled.scala 40:37]
  wire  _GEN_145; // @[HandShaking.scala 716:29]
  wire  _T_75; // @[Decoupled.scala 40:37]
  wire  _GEN_147; // @[HandShaking.scala 716:29]
  wire  _T_76; // @[Decoupled.scala 40:37]
  wire  _GEN_149; // @[HandShaking.scala 716:29]
  wire  _T_77; // @[Decoupled.scala 40:37]
  wire  _GEN_151; // @[HandShaking.scala 716:29]
  wire  _T_78; // @[Decoupled.scala 40:37]
  wire  _GEN_153; // @[HandShaking.scala 716:29]
  wire  _T_79; // @[Decoupled.scala 40:37]
  wire  _GEN_155; // @[HandShaking.scala 716:29]
  wire  _T_80; // @[Decoupled.scala 40:37]
  wire  _GEN_157; // @[HandShaking.scala 716:29]
  wire  _T_81; // @[Decoupled.scala 40:37]
  wire  _GEN_159; // @[HandShaking.scala 716:29]
  wire  _T_82; // @[Decoupled.scala 40:37]
  wire  _GEN_161; // @[HandShaking.scala 716:29]
  wire  _T_83; // @[Decoupled.scala 40:37]
  wire  _GEN_163; // @[HandShaking.scala 716:29]
  wire  _T_84; // @[Decoupled.scala 40:37]
  wire  _GEN_165; // @[HandShaking.scala 716:29]
  wire  _T_85; // @[Decoupled.scala 40:37]
  wire  _GEN_167; // @[HandShaking.scala 716:29]
  wire  _T_86; // @[Decoupled.scala 40:37]
  wire  _GEN_169; // @[HandShaking.scala 716:29]
  wire  _T_87; // @[Decoupled.scala 40:37]
  wire  _GEN_171; // @[HandShaking.scala 716:29]
  wire  _T_88; // @[Decoupled.scala 40:37]
  wire  _GEN_173; // @[HandShaking.scala 716:29]
  wire  _T_89; // @[Decoupled.scala 40:37]
  wire  _GEN_175; // @[HandShaking.scala 716:29]
  wire  _T_90; // @[Decoupled.scala 40:37]
  wire  _GEN_177; // @[HandShaking.scala 716:29]
  wire  _T_91; // @[Decoupled.scala 40:37]
  wire  _GEN_179; // @[HandShaking.scala 716:29]
  wire  _T_92; // @[Decoupled.scala 40:37]
  wire  _GEN_181; // @[HandShaking.scala 716:29]
  wire  _T_93; // @[Decoupled.scala 40:37]
  wire  _GEN_183; // @[HandShaking.scala 716:29]
  wire  _T_94; // @[Decoupled.scala 40:37]
  wire  _GEN_185; // @[HandShaking.scala 716:29]
  wire  _T_95; // @[Decoupled.scala 40:37]
  wire  _GEN_187; // @[HandShaking.scala 727:32]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_187;
  wire [14:0] _T_98; // @[Counter.scala 38:22]
  reg [4:0] predicate_in_R_0_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_188;
  reg  predicate_in_R_0_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_189;
  reg [4:0] predicate_in_R_1_taskID; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_190;
  reg  predicate_in_R_1_control; // @[BasicBlock.scala 64:51]
  reg [31:0] _RAND_191;
  reg  predicate_control_R_0; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_192;
  reg  predicate_control_R_1; // @[BasicBlock.scala 65:36]
  reg [31:0] _RAND_193;
  reg  predicate_valid_R_0; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_194;
  reg  predicate_valid_R_1; // @[BasicBlock.scala 66:54]
  reg [31:0] _RAND_195;
  reg  state; // @[BasicBlock.scala 69:22]
  reg [31:0] _RAND_196;
  wire  predicate; // @[BasicBlock.scala 75:58]
  wire [4:0] predicate_task; // @[BasicBlock.scala 76:62]
  wire  _T_103; // @[Decoupled.scala 40:37]
  wire  _T_104; // @[Decoupled.scala 40:37]
  wire  _T_105; // @[BasicBlock.scala 78:91]
  wire  _T_106; // @[BasicBlock.scala 78:91]
  wire  start; // @[BasicBlock.scala 78:107]
  wire [1:0] _T_111; // @[BasicBlock.scala 102:52]
  wire  _T_112; // @[Conditional.scala 37:30]
  wire  _GEN_197; // @[BasicBlock.scala 112:19]
  wire  _GEN_198; // @[BasicBlock.scala 112:19]
  wire  _GEN_199; // @[BasicBlock.scala 112:19]
  wire  _GEN_200; // @[BasicBlock.scala 112:19]
  wire  _GEN_201; // @[BasicBlock.scala 112:19]
  wire  _GEN_202; // @[BasicBlock.scala 112:19]
  wire  _GEN_203; // @[BasicBlock.scala 112:19]
  wire  _GEN_204; // @[BasicBlock.scala 112:19]
  wire  _GEN_205; // @[BasicBlock.scala 112:19]
  wire  _GEN_206; // @[BasicBlock.scala 112:19]
  wire  _GEN_207; // @[BasicBlock.scala 112:19]
  wire  _GEN_208; // @[BasicBlock.scala 112:19]
  wire  _GEN_209; // @[BasicBlock.scala 112:19]
  wire  _GEN_210; // @[BasicBlock.scala 112:19]
  wire  _GEN_211; // @[BasicBlock.scala 112:19]
  wire  _GEN_212; // @[BasicBlock.scala 112:19]
  wire  _GEN_213; // @[BasicBlock.scala 112:19]
  wire  _GEN_214; // @[BasicBlock.scala 112:19]
  wire  _GEN_215; // @[BasicBlock.scala 112:19]
  wire  _GEN_216; // @[BasicBlock.scala 112:19]
  wire  _GEN_217; // @[BasicBlock.scala 112:19]
  wire  _GEN_218; // @[BasicBlock.scala 112:19]
  wire  _GEN_219; // @[BasicBlock.scala 112:19]
  wire  _GEN_220; // @[BasicBlock.scala 112:19]
  wire  _GEN_221; // @[BasicBlock.scala 112:19]
  wire  _GEN_222; // @[BasicBlock.scala 112:19]
  wire  _GEN_223; // @[BasicBlock.scala 112:19]
  wire  _GEN_224; // @[BasicBlock.scala 112:19]
  wire  _GEN_225; // @[BasicBlock.scala 112:19]
  wire  _GEN_226; // @[BasicBlock.scala 112:19]
  wire  _GEN_227; // @[BasicBlock.scala 112:19]
  wire  _GEN_228; // @[BasicBlock.scala 112:19]
  wire  _GEN_229; // @[BasicBlock.scala 112:19]
  wire  _GEN_230; // @[BasicBlock.scala 112:19]
  wire  _GEN_231; // @[BasicBlock.scala 112:19]
  wire  _GEN_232; // @[BasicBlock.scala 112:19]
  wire  _GEN_233; // @[BasicBlock.scala 112:19]
  wire  _GEN_234; // @[BasicBlock.scala 112:19]
  wire  _GEN_235; // @[BasicBlock.scala 112:19]
  wire  _GEN_236; // @[BasicBlock.scala 112:19]
  wire  _GEN_237; // @[BasicBlock.scala 112:19]
  wire  _GEN_238; // @[BasicBlock.scala 112:19]
  wire  _GEN_239; // @[BasicBlock.scala 112:19]
  wire  _GEN_240; // @[BasicBlock.scala 112:19]
  wire  _GEN_241; // @[BasicBlock.scala 112:19]
  wire  _GEN_242; // @[BasicBlock.scala 112:19]
  wire  _GEN_243; // @[BasicBlock.scala 112:19]
  wire  _GEN_244; // @[BasicBlock.scala 112:19]
  wire  _GEN_245; // @[BasicBlock.scala 112:19]
  wire  _GEN_246; // @[BasicBlock.scala 112:19]
  wire  _GEN_247; // @[BasicBlock.scala 112:19]
  wire  _GEN_248; // @[BasicBlock.scala 112:19]
  wire  _GEN_249; // @[BasicBlock.scala 112:19]
  wire  _GEN_250; // @[BasicBlock.scala 112:19]
  wire  _GEN_251; // @[BasicBlock.scala 112:19]
  wire  _GEN_252; // @[BasicBlock.scala 112:19]
  wire  _GEN_253; // @[BasicBlock.scala 112:19]
  wire  _GEN_254; // @[BasicBlock.scala 112:19]
  wire  _GEN_255; // @[BasicBlock.scala 112:19]
  wire  _GEN_256; // @[BasicBlock.scala 112:19]
  wire  _GEN_257; // @[BasicBlock.scala 112:19]
  wire  _GEN_258; // @[BasicBlock.scala 112:19]
  wire  _GEN_259; // @[BasicBlock.scala 112:19]
  wire  _GEN_260; // @[BasicBlock.scala 112:19]
  wire  _GEN_261; // @[BasicBlock.scala 112:19]
  wire  _GEN_262; // @[BasicBlock.scala 112:19]
  wire  _GEN_263; // @[BasicBlock.scala 112:19]
  wire  _GEN_264; // @[BasicBlock.scala 112:19]
  wire  _GEN_265; // @[BasicBlock.scala 112:19]
  wire  _GEN_266; // @[BasicBlock.scala 112:19]
  wire  _GEN_267; // @[BasicBlock.scala 112:19]
  wire  _GEN_268; // @[BasicBlock.scala 112:19]
  wire  _GEN_269; // @[BasicBlock.scala 112:19]
  wire  _GEN_270; // @[BasicBlock.scala 112:19]
  wire  _GEN_271; // @[BasicBlock.scala 112:19]
  wire  _GEN_272; // @[BasicBlock.scala 112:19]
  wire  _GEN_273; // @[BasicBlock.scala 112:19]
  wire  _GEN_274; // @[BasicBlock.scala 112:19]
  wire  _GEN_275; // @[BasicBlock.scala 112:19]
  wire  _GEN_276; // @[BasicBlock.scala 112:19]
  wire  _GEN_277; // @[BasicBlock.scala 112:19]
  wire  _GEN_278; // @[BasicBlock.scala 112:19]
  wire  _GEN_279; // @[BasicBlock.scala 112:19]
  wire  _GEN_280; // @[BasicBlock.scala 112:19]
  wire  _GEN_281; // @[BasicBlock.scala 112:19]
  wire  _GEN_282; // @[BasicBlock.scala 112:19]
  wire  _GEN_283; // @[BasicBlock.scala 112:19]
  wire  _GEN_284; // @[BasicBlock.scala 112:19]
  wire  _GEN_285; // @[BasicBlock.scala 112:19]
  wire  _GEN_286; // @[BasicBlock.scala 112:19]
  wire  _GEN_287; // @[BasicBlock.scala 112:19]
  wire  _GEN_288; // @[BasicBlock.scala 112:19]
  wire  _GEN_289; // @[BasicBlock.scala 112:19]
  wire  _GEN_290; // @[BasicBlock.scala 112:19]
  wire  _GEN_291; // @[BasicBlock.scala 112:19]
  wire [4:0] _T_118; // @[HandShaking.scala 741:17]
  wire [10:0] _T_124; // @[HandShaking.scala 741:17]
  wire [5:0] _T_129; // @[HandShaking.scala 741:17]
  wire [22:0] _T_136; // @[HandShaking.scala 741:17]
  wire [4:0] _T_140; // @[HandShaking.scala 741:17]
  wire [10:0] _T_146; // @[HandShaking.scala 741:17]
  wire [5:0] _T_151; // @[HandShaking.scala 741:17]
  wire [45:0] _T_159; // @[HandShaking.scala 741:17]
  wire [4:0] _T_163; // @[HandShaking.scala 741:17]
  wire [10:0] _T_169; // @[HandShaking.scala 741:17]
  wire [5:0] _T_174; // @[HandShaking.scala 741:17]
  wire [22:0] _T_181; // @[HandShaking.scala 741:17]
  wire [5:0] _T_186; // @[HandShaking.scala 741:17]
  wire [11:0] _T_192; // @[HandShaking.scala 741:17]
  wire [5:0] _T_197; // @[HandShaking.scala 741:17]
  wire [92:0] _T_206; // @[HandShaking.scala 741:17]
  wire  _T_207; // @[HandShaking.scala 741:24]
  wire  _T_210; // @[BasicBlock.scala 126:19]
  wire  _T_211; // @[BasicBlock.scala 126:19]
  wire  _GEN_677; // @[BasicBlock.scala 126:19]
  wire  _GEN_678; // @[BasicBlock.scala 126:19]
  wire  _GEN_679; // @[BasicBlock.scala 126:19]
  wire  _GEN_680; // @[BasicBlock.scala 126:19]
  wire  _GEN_684; // @[BasicBlock.scala 132:19]
  wire  _GEN_685; // @[BasicBlock.scala 132:19]
  assign _T_2 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_1 = _T_2 ? 1'h0 : out_valid_R_0; // @[HandShaking.scala 716:29]
  assign _T_3 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_3 = _T_3 ? 1'h0 : out_valid_R_1; // @[HandShaking.scala 716:29]
  assign _T_4 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_4 ? 1'h0 : out_valid_R_2; // @[HandShaking.scala 716:29]
  assign _T_5 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_5 ? 1'h0 : out_valid_R_3; // @[HandShaking.scala 716:29]
  assign _T_6 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_6 ? 1'h0 : out_valid_R_4; // @[HandShaking.scala 716:29]
  assign _T_7 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_7 ? 1'h0 : out_valid_R_5; // @[HandShaking.scala 716:29]
  assign _T_8 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_8 ? 1'h0 : out_valid_R_6; // @[HandShaking.scala 716:29]
  assign _T_9 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_9 ? 1'h0 : out_valid_R_7; // @[HandShaking.scala 716:29]
  assign _T_10 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_10 ? 1'h0 : out_valid_R_8; // @[HandShaking.scala 716:29]
  assign _T_11 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_11 ? 1'h0 : out_valid_R_9; // @[HandShaking.scala 716:29]
  assign _T_12 = io_Out_10_ready & io_Out_10_valid; // @[Decoupled.scala 40:37]
  assign _GEN_21 = _T_12 ? 1'h0 : out_valid_R_10; // @[HandShaking.scala 716:29]
  assign _T_13 = io_Out_11_ready & io_Out_11_valid; // @[Decoupled.scala 40:37]
  assign _GEN_23 = _T_13 ? 1'h0 : out_valid_R_11; // @[HandShaking.scala 716:29]
  assign _T_14 = io_Out_12_ready & io_Out_12_valid; // @[Decoupled.scala 40:37]
  assign _GEN_25 = _T_14 ? 1'h0 : out_valid_R_12; // @[HandShaking.scala 716:29]
  assign _T_15 = io_Out_13_ready & io_Out_13_valid; // @[Decoupled.scala 40:37]
  assign _GEN_27 = _T_15 ? 1'h0 : out_valid_R_13; // @[HandShaking.scala 716:29]
  assign _T_16 = io_Out_14_ready & io_Out_14_valid; // @[Decoupled.scala 40:37]
  assign _GEN_29 = _T_16 ? 1'h0 : out_valid_R_14; // @[HandShaking.scala 716:29]
  assign _T_17 = io_Out_15_ready & io_Out_15_valid; // @[Decoupled.scala 40:37]
  assign _GEN_31 = _T_17 ? 1'h0 : out_valid_R_15; // @[HandShaking.scala 716:29]
  assign _T_18 = io_Out_16_ready & io_Out_16_valid; // @[Decoupled.scala 40:37]
  assign _GEN_33 = _T_18 ? 1'h0 : out_valid_R_16; // @[HandShaking.scala 716:29]
  assign _T_19 = io_Out_17_ready & io_Out_17_valid; // @[Decoupled.scala 40:37]
  assign _GEN_35 = _T_19 ? 1'h0 : out_valid_R_17; // @[HandShaking.scala 716:29]
  assign _T_20 = io_Out_18_ready & io_Out_18_valid; // @[Decoupled.scala 40:37]
  assign _GEN_37 = _T_20 ? 1'h0 : out_valid_R_18; // @[HandShaking.scala 716:29]
  assign _T_21 = io_Out_19_ready & io_Out_19_valid; // @[Decoupled.scala 40:37]
  assign _GEN_39 = _T_21 ? 1'h0 : out_valid_R_19; // @[HandShaking.scala 716:29]
  assign _T_22 = io_Out_20_ready & io_Out_20_valid; // @[Decoupled.scala 40:37]
  assign _GEN_41 = _T_22 ? 1'h0 : out_valid_R_20; // @[HandShaking.scala 716:29]
  assign _T_23 = io_Out_21_ready & io_Out_21_valid; // @[Decoupled.scala 40:37]
  assign _GEN_43 = _T_23 ? 1'h0 : out_valid_R_21; // @[HandShaking.scala 716:29]
  assign _T_24 = io_Out_22_ready & io_Out_22_valid; // @[Decoupled.scala 40:37]
  assign _GEN_45 = _T_24 ? 1'h0 : out_valid_R_22; // @[HandShaking.scala 716:29]
  assign _T_25 = io_Out_23_ready & io_Out_23_valid; // @[Decoupled.scala 40:37]
  assign _GEN_47 = _T_25 ? 1'h0 : out_valid_R_23; // @[HandShaking.scala 716:29]
  assign _T_26 = io_Out_24_ready & io_Out_24_valid; // @[Decoupled.scala 40:37]
  assign _GEN_49 = _T_26 ? 1'h0 : out_valid_R_24; // @[HandShaking.scala 716:29]
  assign _T_27 = io_Out_25_ready & io_Out_25_valid; // @[Decoupled.scala 40:37]
  assign _GEN_51 = _T_27 ? 1'h0 : out_valid_R_25; // @[HandShaking.scala 716:29]
  assign _T_28 = io_Out_26_ready & io_Out_26_valid; // @[Decoupled.scala 40:37]
  assign _GEN_53 = _T_28 ? 1'h0 : out_valid_R_26; // @[HandShaking.scala 716:29]
  assign _T_29 = io_Out_27_ready & io_Out_27_valid; // @[Decoupled.scala 40:37]
  assign _GEN_55 = _T_29 ? 1'h0 : out_valid_R_27; // @[HandShaking.scala 716:29]
  assign _T_30 = io_Out_28_ready & io_Out_28_valid; // @[Decoupled.scala 40:37]
  assign _GEN_57 = _T_30 ? 1'h0 : out_valid_R_28; // @[HandShaking.scala 716:29]
  assign _T_31 = io_Out_29_ready & io_Out_29_valid; // @[Decoupled.scala 40:37]
  assign _GEN_59 = _T_31 ? 1'h0 : out_valid_R_29; // @[HandShaking.scala 716:29]
  assign _T_32 = io_Out_30_ready & io_Out_30_valid; // @[Decoupled.scala 40:37]
  assign _GEN_61 = _T_32 ? 1'h0 : out_valid_R_30; // @[HandShaking.scala 716:29]
  assign _T_33 = io_Out_31_ready & io_Out_31_valid; // @[Decoupled.scala 40:37]
  assign _GEN_63 = _T_33 ? 1'h0 : out_valid_R_31; // @[HandShaking.scala 716:29]
  assign _T_34 = io_Out_32_ready & io_Out_32_valid; // @[Decoupled.scala 40:37]
  assign _GEN_65 = _T_34 ? 1'h0 : out_valid_R_32; // @[HandShaking.scala 716:29]
  assign _T_35 = io_Out_33_ready & io_Out_33_valid; // @[Decoupled.scala 40:37]
  assign _GEN_67 = _T_35 ? 1'h0 : out_valid_R_33; // @[HandShaking.scala 716:29]
  assign _T_36 = io_Out_34_ready & io_Out_34_valid; // @[Decoupled.scala 40:37]
  assign _GEN_69 = _T_36 ? 1'h0 : out_valid_R_34; // @[HandShaking.scala 716:29]
  assign _T_37 = io_Out_35_ready & io_Out_35_valid; // @[Decoupled.scala 40:37]
  assign _GEN_71 = _T_37 ? 1'h0 : out_valid_R_35; // @[HandShaking.scala 716:29]
  assign _T_38 = io_Out_36_ready & io_Out_36_valid; // @[Decoupled.scala 40:37]
  assign _GEN_73 = _T_38 ? 1'h0 : out_valid_R_36; // @[HandShaking.scala 716:29]
  assign _T_39 = io_Out_37_ready & io_Out_37_valid; // @[Decoupled.scala 40:37]
  assign _GEN_75 = _T_39 ? 1'h0 : out_valid_R_37; // @[HandShaking.scala 716:29]
  assign _T_40 = io_Out_38_ready & io_Out_38_valid; // @[Decoupled.scala 40:37]
  assign _GEN_77 = _T_40 ? 1'h0 : out_valid_R_38; // @[HandShaking.scala 716:29]
  assign _T_41 = io_Out_39_ready & io_Out_39_valid; // @[Decoupled.scala 40:37]
  assign _GEN_79 = _T_41 ? 1'h0 : out_valid_R_39; // @[HandShaking.scala 716:29]
  assign _T_42 = io_Out_40_ready & io_Out_40_valid; // @[Decoupled.scala 40:37]
  assign _GEN_81 = _T_42 ? 1'h0 : out_valid_R_40; // @[HandShaking.scala 716:29]
  assign _T_43 = io_Out_41_ready & io_Out_41_valid; // @[Decoupled.scala 40:37]
  assign _GEN_83 = _T_43 ? 1'h0 : out_valid_R_41; // @[HandShaking.scala 716:29]
  assign _T_44 = io_Out_42_ready & io_Out_42_valid; // @[Decoupled.scala 40:37]
  assign _GEN_85 = _T_44 ? 1'h0 : out_valid_R_42; // @[HandShaking.scala 716:29]
  assign _T_45 = io_Out_43_ready & io_Out_43_valid; // @[Decoupled.scala 40:37]
  assign _GEN_87 = _T_45 ? 1'h0 : out_valid_R_43; // @[HandShaking.scala 716:29]
  assign _T_46 = io_Out_44_ready & io_Out_44_valid; // @[Decoupled.scala 40:37]
  assign _GEN_89 = _T_46 ? 1'h0 : out_valid_R_44; // @[HandShaking.scala 716:29]
  assign _T_47 = io_Out_45_ready & io_Out_45_valid; // @[Decoupled.scala 40:37]
  assign _GEN_91 = _T_47 ? 1'h0 : out_valid_R_45; // @[HandShaking.scala 716:29]
  assign _T_48 = io_Out_46_ready & io_Out_46_valid; // @[Decoupled.scala 40:37]
  assign _GEN_93 = _T_48 ? 1'h0 : out_valid_R_46; // @[HandShaking.scala 716:29]
  assign _T_49 = io_Out_47_ready & io_Out_47_valid; // @[Decoupled.scala 40:37]
  assign _GEN_95 = _T_49 ? 1'h0 : out_valid_R_47; // @[HandShaking.scala 716:29]
  assign _T_50 = io_Out_48_ready & io_Out_48_valid; // @[Decoupled.scala 40:37]
  assign _GEN_97 = _T_50 ? 1'h0 : out_valid_R_48; // @[HandShaking.scala 716:29]
  assign _T_51 = io_Out_49_ready & io_Out_49_valid; // @[Decoupled.scala 40:37]
  assign _GEN_99 = _T_51 ? 1'h0 : out_valid_R_49; // @[HandShaking.scala 716:29]
  assign _T_52 = io_Out_50_ready & io_Out_50_valid; // @[Decoupled.scala 40:37]
  assign _GEN_101 = _T_52 ? 1'h0 : out_valid_R_50; // @[HandShaking.scala 716:29]
  assign _T_53 = io_Out_51_ready & io_Out_51_valid; // @[Decoupled.scala 40:37]
  assign _GEN_103 = _T_53 ? 1'h0 : out_valid_R_51; // @[HandShaking.scala 716:29]
  assign _T_54 = io_Out_52_ready & io_Out_52_valid; // @[Decoupled.scala 40:37]
  assign _GEN_105 = _T_54 ? 1'h0 : out_valid_R_52; // @[HandShaking.scala 716:29]
  assign _T_55 = io_Out_53_ready & io_Out_53_valid; // @[Decoupled.scala 40:37]
  assign _GEN_107 = _T_55 ? 1'h0 : out_valid_R_53; // @[HandShaking.scala 716:29]
  assign _T_56 = io_Out_54_ready & io_Out_54_valid; // @[Decoupled.scala 40:37]
  assign _GEN_109 = _T_56 ? 1'h0 : out_valid_R_54; // @[HandShaking.scala 716:29]
  assign _T_57 = io_Out_55_ready & io_Out_55_valid; // @[Decoupled.scala 40:37]
  assign _GEN_111 = _T_57 ? 1'h0 : out_valid_R_55; // @[HandShaking.scala 716:29]
  assign _T_58 = io_Out_56_ready & io_Out_56_valid; // @[Decoupled.scala 40:37]
  assign _GEN_113 = _T_58 ? 1'h0 : out_valid_R_56; // @[HandShaking.scala 716:29]
  assign _T_59 = io_Out_57_ready & io_Out_57_valid; // @[Decoupled.scala 40:37]
  assign _GEN_115 = _T_59 ? 1'h0 : out_valid_R_57; // @[HandShaking.scala 716:29]
  assign _T_60 = io_Out_58_ready & io_Out_58_valid; // @[Decoupled.scala 40:37]
  assign _GEN_117 = _T_60 ? 1'h0 : out_valid_R_58; // @[HandShaking.scala 716:29]
  assign _T_61 = io_Out_59_ready & io_Out_59_valid; // @[Decoupled.scala 40:37]
  assign _GEN_119 = _T_61 ? 1'h0 : out_valid_R_59; // @[HandShaking.scala 716:29]
  assign _T_62 = io_Out_60_ready & io_Out_60_valid; // @[Decoupled.scala 40:37]
  assign _GEN_121 = _T_62 ? 1'h0 : out_valid_R_60; // @[HandShaking.scala 716:29]
  assign _T_63 = io_Out_61_ready & io_Out_61_valid; // @[Decoupled.scala 40:37]
  assign _GEN_123 = _T_63 ? 1'h0 : out_valid_R_61; // @[HandShaking.scala 716:29]
  assign _T_64 = io_Out_62_ready & io_Out_62_valid; // @[Decoupled.scala 40:37]
  assign _GEN_125 = _T_64 ? 1'h0 : out_valid_R_62; // @[HandShaking.scala 716:29]
  assign _T_65 = io_Out_63_ready & io_Out_63_valid; // @[Decoupled.scala 40:37]
  assign _GEN_127 = _T_65 ? 1'h0 : out_valid_R_63; // @[HandShaking.scala 716:29]
  assign _T_66 = io_Out_64_ready & io_Out_64_valid; // @[Decoupled.scala 40:37]
  assign _GEN_129 = _T_66 ? 1'h0 : out_valid_R_64; // @[HandShaking.scala 716:29]
  assign _T_67 = io_Out_65_ready & io_Out_65_valid; // @[Decoupled.scala 40:37]
  assign _GEN_131 = _T_67 ? 1'h0 : out_valid_R_65; // @[HandShaking.scala 716:29]
  assign _T_68 = io_Out_66_ready & io_Out_66_valid; // @[Decoupled.scala 40:37]
  assign _GEN_133 = _T_68 ? 1'h0 : out_valid_R_66; // @[HandShaking.scala 716:29]
  assign _T_69 = io_Out_67_ready & io_Out_67_valid; // @[Decoupled.scala 40:37]
  assign _GEN_135 = _T_69 ? 1'h0 : out_valid_R_67; // @[HandShaking.scala 716:29]
  assign _T_70 = io_Out_68_ready & io_Out_68_valid; // @[Decoupled.scala 40:37]
  assign _GEN_137 = _T_70 ? 1'h0 : out_valid_R_68; // @[HandShaking.scala 716:29]
  assign _T_71 = io_Out_69_ready & io_Out_69_valid; // @[Decoupled.scala 40:37]
  assign _GEN_139 = _T_71 ? 1'h0 : out_valid_R_69; // @[HandShaking.scala 716:29]
  assign _T_72 = io_Out_70_ready & io_Out_70_valid; // @[Decoupled.scala 40:37]
  assign _GEN_141 = _T_72 ? 1'h0 : out_valid_R_70; // @[HandShaking.scala 716:29]
  assign _T_73 = io_Out_71_ready & io_Out_71_valid; // @[Decoupled.scala 40:37]
  assign _GEN_143 = _T_73 ? 1'h0 : out_valid_R_71; // @[HandShaking.scala 716:29]
  assign _T_74 = io_Out_72_ready & io_Out_72_valid; // @[Decoupled.scala 40:37]
  assign _GEN_145 = _T_74 ? 1'h0 : out_valid_R_72; // @[HandShaking.scala 716:29]
  assign _T_75 = io_Out_73_ready & io_Out_73_valid; // @[Decoupled.scala 40:37]
  assign _GEN_147 = _T_75 ? 1'h0 : out_valid_R_73; // @[HandShaking.scala 716:29]
  assign _T_76 = io_Out_74_ready & io_Out_74_valid; // @[Decoupled.scala 40:37]
  assign _GEN_149 = _T_76 ? 1'h0 : out_valid_R_74; // @[HandShaking.scala 716:29]
  assign _T_77 = io_Out_75_ready & io_Out_75_valid; // @[Decoupled.scala 40:37]
  assign _GEN_151 = _T_77 ? 1'h0 : out_valid_R_75; // @[HandShaking.scala 716:29]
  assign _T_78 = io_Out_76_ready & io_Out_76_valid; // @[Decoupled.scala 40:37]
  assign _GEN_153 = _T_78 ? 1'h0 : out_valid_R_76; // @[HandShaking.scala 716:29]
  assign _T_79 = io_Out_77_ready & io_Out_77_valid; // @[Decoupled.scala 40:37]
  assign _GEN_155 = _T_79 ? 1'h0 : out_valid_R_77; // @[HandShaking.scala 716:29]
  assign _T_80 = io_Out_78_ready & io_Out_78_valid; // @[Decoupled.scala 40:37]
  assign _GEN_157 = _T_80 ? 1'h0 : out_valid_R_78; // @[HandShaking.scala 716:29]
  assign _T_81 = io_Out_79_ready & io_Out_79_valid; // @[Decoupled.scala 40:37]
  assign _GEN_159 = _T_81 ? 1'h0 : out_valid_R_79; // @[HandShaking.scala 716:29]
  assign _T_82 = io_Out_80_ready & io_Out_80_valid; // @[Decoupled.scala 40:37]
  assign _GEN_161 = _T_82 ? 1'h0 : out_valid_R_80; // @[HandShaking.scala 716:29]
  assign _T_83 = io_Out_81_ready & io_Out_81_valid; // @[Decoupled.scala 40:37]
  assign _GEN_163 = _T_83 ? 1'h0 : out_valid_R_81; // @[HandShaking.scala 716:29]
  assign _T_84 = io_Out_82_ready & io_Out_82_valid; // @[Decoupled.scala 40:37]
  assign _GEN_165 = _T_84 ? 1'h0 : out_valid_R_82; // @[HandShaking.scala 716:29]
  assign _T_85 = io_Out_83_ready & io_Out_83_valid; // @[Decoupled.scala 40:37]
  assign _GEN_167 = _T_85 ? 1'h0 : out_valid_R_83; // @[HandShaking.scala 716:29]
  assign _T_86 = io_Out_84_ready & io_Out_84_valid; // @[Decoupled.scala 40:37]
  assign _GEN_169 = _T_86 ? 1'h0 : out_valid_R_84; // @[HandShaking.scala 716:29]
  assign _T_87 = io_Out_85_ready & io_Out_85_valid; // @[Decoupled.scala 40:37]
  assign _GEN_171 = _T_87 ? 1'h0 : out_valid_R_85; // @[HandShaking.scala 716:29]
  assign _T_88 = io_Out_86_ready & io_Out_86_valid; // @[Decoupled.scala 40:37]
  assign _GEN_173 = _T_88 ? 1'h0 : out_valid_R_86; // @[HandShaking.scala 716:29]
  assign _T_89 = io_Out_87_ready & io_Out_87_valid; // @[Decoupled.scala 40:37]
  assign _GEN_175 = _T_89 ? 1'h0 : out_valid_R_87; // @[HandShaking.scala 716:29]
  assign _T_90 = io_Out_88_ready & io_Out_88_valid; // @[Decoupled.scala 40:37]
  assign _GEN_177 = _T_90 ? 1'h0 : out_valid_R_88; // @[HandShaking.scala 716:29]
  assign _T_91 = io_Out_89_ready & io_Out_89_valid; // @[Decoupled.scala 40:37]
  assign _GEN_179 = _T_91 ? 1'h0 : out_valid_R_89; // @[HandShaking.scala 716:29]
  assign _T_92 = io_Out_90_ready & io_Out_90_valid; // @[Decoupled.scala 40:37]
  assign _GEN_181 = _T_92 ? 1'h0 : out_valid_R_90; // @[HandShaking.scala 716:29]
  assign _T_93 = io_Out_91_ready & io_Out_91_valid; // @[Decoupled.scala 40:37]
  assign _GEN_183 = _T_93 ? 1'h0 : out_valid_R_91; // @[HandShaking.scala 716:29]
  assign _T_94 = io_Out_92_ready & io_Out_92_valid; // @[Decoupled.scala 40:37]
  assign _GEN_185 = _T_94 ? 1'h0 : out_valid_R_92; // @[HandShaking.scala 716:29]
  assign _T_95 = io_MaskBB_0_ready & io_MaskBB_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_187 = _T_95 ? 1'h0 : mask_valid_R_0; // @[HandShaking.scala 727:32]
  assign _T_98 = value + 15'h1; // @[Counter.scala 38:22]
  assign predicate = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 75:58]
  assign predicate_task = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 76:62]
  assign _T_103 = io_predicateIn_0_ready & io_predicateIn_0_valid; // @[Decoupled.scala 40:37]
  assign _T_104 = io_predicateIn_1_ready & io_predicateIn_1_valid; // @[Decoupled.scala 40:37]
  assign _T_105 = _T_103 | predicate_valid_R_0; // @[BasicBlock.scala 78:91]
  assign _T_106 = _T_104 | predicate_valid_R_1; // @[BasicBlock.scala 78:91]
  assign start = _T_105 & _T_106; // @[BasicBlock.scala 78:107]
  assign _T_111 = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:52]
  assign _T_112 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_197 = start | _GEN_1; // @[BasicBlock.scala 112:19]
  assign _GEN_198 = start | _GEN_3; // @[BasicBlock.scala 112:19]
  assign _GEN_199 = start | _GEN_5; // @[BasicBlock.scala 112:19]
  assign _GEN_200 = start | _GEN_7; // @[BasicBlock.scala 112:19]
  assign _GEN_201 = start | _GEN_9; // @[BasicBlock.scala 112:19]
  assign _GEN_202 = start | _GEN_11; // @[BasicBlock.scala 112:19]
  assign _GEN_203 = start | _GEN_13; // @[BasicBlock.scala 112:19]
  assign _GEN_204 = start | _GEN_15; // @[BasicBlock.scala 112:19]
  assign _GEN_205 = start | _GEN_17; // @[BasicBlock.scala 112:19]
  assign _GEN_206 = start | _GEN_19; // @[BasicBlock.scala 112:19]
  assign _GEN_207 = start | _GEN_21; // @[BasicBlock.scala 112:19]
  assign _GEN_208 = start | _GEN_23; // @[BasicBlock.scala 112:19]
  assign _GEN_209 = start | _GEN_25; // @[BasicBlock.scala 112:19]
  assign _GEN_210 = start | _GEN_27; // @[BasicBlock.scala 112:19]
  assign _GEN_211 = start | _GEN_29; // @[BasicBlock.scala 112:19]
  assign _GEN_212 = start | _GEN_31; // @[BasicBlock.scala 112:19]
  assign _GEN_213 = start | _GEN_33; // @[BasicBlock.scala 112:19]
  assign _GEN_214 = start | _GEN_35; // @[BasicBlock.scala 112:19]
  assign _GEN_215 = start | _GEN_37; // @[BasicBlock.scala 112:19]
  assign _GEN_216 = start | _GEN_39; // @[BasicBlock.scala 112:19]
  assign _GEN_217 = start | _GEN_41; // @[BasicBlock.scala 112:19]
  assign _GEN_218 = start | _GEN_43; // @[BasicBlock.scala 112:19]
  assign _GEN_219 = start | _GEN_45; // @[BasicBlock.scala 112:19]
  assign _GEN_220 = start | _GEN_47; // @[BasicBlock.scala 112:19]
  assign _GEN_221 = start | _GEN_49; // @[BasicBlock.scala 112:19]
  assign _GEN_222 = start | _GEN_51; // @[BasicBlock.scala 112:19]
  assign _GEN_223 = start | _GEN_53; // @[BasicBlock.scala 112:19]
  assign _GEN_224 = start | _GEN_55; // @[BasicBlock.scala 112:19]
  assign _GEN_225 = start | _GEN_57; // @[BasicBlock.scala 112:19]
  assign _GEN_226 = start | _GEN_59; // @[BasicBlock.scala 112:19]
  assign _GEN_227 = start | _GEN_61; // @[BasicBlock.scala 112:19]
  assign _GEN_228 = start | _GEN_63; // @[BasicBlock.scala 112:19]
  assign _GEN_229 = start | _GEN_65; // @[BasicBlock.scala 112:19]
  assign _GEN_230 = start | _GEN_67; // @[BasicBlock.scala 112:19]
  assign _GEN_231 = start | _GEN_69; // @[BasicBlock.scala 112:19]
  assign _GEN_232 = start | _GEN_71; // @[BasicBlock.scala 112:19]
  assign _GEN_233 = start | _GEN_73; // @[BasicBlock.scala 112:19]
  assign _GEN_234 = start | _GEN_75; // @[BasicBlock.scala 112:19]
  assign _GEN_235 = start | _GEN_77; // @[BasicBlock.scala 112:19]
  assign _GEN_236 = start | _GEN_79; // @[BasicBlock.scala 112:19]
  assign _GEN_237 = start | _GEN_81; // @[BasicBlock.scala 112:19]
  assign _GEN_238 = start | _GEN_83; // @[BasicBlock.scala 112:19]
  assign _GEN_239 = start | _GEN_85; // @[BasicBlock.scala 112:19]
  assign _GEN_240 = start | _GEN_87; // @[BasicBlock.scala 112:19]
  assign _GEN_241 = start | _GEN_89; // @[BasicBlock.scala 112:19]
  assign _GEN_242 = start | _GEN_91; // @[BasicBlock.scala 112:19]
  assign _GEN_243 = start | _GEN_93; // @[BasicBlock.scala 112:19]
  assign _GEN_244 = start | _GEN_95; // @[BasicBlock.scala 112:19]
  assign _GEN_245 = start | _GEN_97; // @[BasicBlock.scala 112:19]
  assign _GEN_246 = start | _GEN_99; // @[BasicBlock.scala 112:19]
  assign _GEN_247 = start | _GEN_101; // @[BasicBlock.scala 112:19]
  assign _GEN_248 = start | _GEN_103; // @[BasicBlock.scala 112:19]
  assign _GEN_249 = start | _GEN_105; // @[BasicBlock.scala 112:19]
  assign _GEN_250 = start | _GEN_107; // @[BasicBlock.scala 112:19]
  assign _GEN_251 = start | _GEN_109; // @[BasicBlock.scala 112:19]
  assign _GEN_252 = start | _GEN_111; // @[BasicBlock.scala 112:19]
  assign _GEN_253 = start | _GEN_113; // @[BasicBlock.scala 112:19]
  assign _GEN_254 = start | _GEN_115; // @[BasicBlock.scala 112:19]
  assign _GEN_255 = start | _GEN_117; // @[BasicBlock.scala 112:19]
  assign _GEN_256 = start | _GEN_119; // @[BasicBlock.scala 112:19]
  assign _GEN_257 = start | _GEN_121; // @[BasicBlock.scala 112:19]
  assign _GEN_258 = start | _GEN_123; // @[BasicBlock.scala 112:19]
  assign _GEN_259 = start | _GEN_125; // @[BasicBlock.scala 112:19]
  assign _GEN_260 = start | _GEN_127; // @[BasicBlock.scala 112:19]
  assign _GEN_261 = start | _GEN_129; // @[BasicBlock.scala 112:19]
  assign _GEN_262 = start | _GEN_131; // @[BasicBlock.scala 112:19]
  assign _GEN_263 = start | _GEN_133; // @[BasicBlock.scala 112:19]
  assign _GEN_264 = start | _GEN_135; // @[BasicBlock.scala 112:19]
  assign _GEN_265 = start | _GEN_137; // @[BasicBlock.scala 112:19]
  assign _GEN_266 = start | _GEN_139; // @[BasicBlock.scala 112:19]
  assign _GEN_267 = start | _GEN_141; // @[BasicBlock.scala 112:19]
  assign _GEN_268 = start | _GEN_143; // @[BasicBlock.scala 112:19]
  assign _GEN_269 = start | _GEN_145; // @[BasicBlock.scala 112:19]
  assign _GEN_270 = start | _GEN_147; // @[BasicBlock.scala 112:19]
  assign _GEN_271 = start | _GEN_149; // @[BasicBlock.scala 112:19]
  assign _GEN_272 = start | _GEN_151; // @[BasicBlock.scala 112:19]
  assign _GEN_273 = start | _GEN_153; // @[BasicBlock.scala 112:19]
  assign _GEN_274 = start | _GEN_155; // @[BasicBlock.scala 112:19]
  assign _GEN_275 = start | _GEN_157; // @[BasicBlock.scala 112:19]
  assign _GEN_276 = start | _GEN_159; // @[BasicBlock.scala 112:19]
  assign _GEN_277 = start | _GEN_161; // @[BasicBlock.scala 112:19]
  assign _GEN_278 = start | _GEN_163; // @[BasicBlock.scala 112:19]
  assign _GEN_279 = start | _GEN_165; // @[BasicBlock.scala 112:19]
  assign _GEN_280 = start | _GEN_167; // @[BasicBlock.scala 112:19]
  assign _GEN_281 = start | _GEN_169; // @[BasicBlock.scala 112:19]
  assign _GEN_282 = start | _GEN_171; // @[BasicBlock.scala 112:19]
  assign _GEN_283 = start | _GEN_173; // @[BasicBlock.scala 112:19]
  assign _GEN_284 = start | _GEN_175; // @[BasicBlock.scala 112:19]
  assign _GEN_285 = start | _GEN_177; // @[BasicBlock.scala 112:19]
  assign _GEN_286 = start | _GEN_179; // @[BasicBlock.scala 112:19]
  assign _GEN_287 = start | _GEN_181; // @[BasicBlock.scala 112:19]
  assign _GEN_288 = start | _GEN_183; // @[BasicBlock.scala 112:19]
  assign _GEN_289 = start | _GEN_185; // @[BasicBlock.scala 112:19]
  assign _GEN_290 = start | _GEN_187; // @[BasicBlock.scala 112:19]
  assign _GEN_291 = start | state; // @[BasicBlock.scala 112:19]
  assign _T_118 = {out_ready_R_4,out_ready_R_3,out_ready_R_2,out_ready_R_1,out_ready_R_0}; // @[HandShaking.scala 741:17]
  assign _T_124 = {out_ready_R_10,out_ready_R_9,out_ready_R_8,out_ready_R_7,out_ready_R_6,out_ready_R_5,_T_118}; // @[HandShaking.scala 741:17]
  assign _T_129 = {out_ready_R_16,out_ready_R_15,out_ready_R_14,out_ready_R_13,out_ready_R_12,out_ready_R_11}; // @[HandShaking.scala 741:17]
  assign _T_136 = {out_ready_R_22,out_ready_R_21,out_ready_R_20,out_ready_R_19,out_ready_R_18,out_ready_R_17,_T_129,_T_124}; // @[HandShaking.scala 741:17]
  assign _T_140 = {out_ready_R_27,out_ready_R_26,out_ready_R_25,out_ready_R_24,out_ready_R_23}; // @[HandShaking.scala 741:17]
  assign _T_146 = {out_ready_R_33,out_ready_R_32,out_ready_R_31,out_ready_R_30,out_ready_R_29,out_ready_R_28,_T_140}; // @[HandShaking.scala 741:17]
  assign _T_151 = {out_ready_R_39,out_ready_R_38,out_ready_R_37,out_ready_R_36,out_ready_R_35,out_ready_R_34}; // @[HandShaking.scala 741:17]
  assign _T_159 = {out_ready_R_45,out_ready_R_44,out_ready_R_43,out_ready_R_42,out_ready_R_41,out_ready_R_40,_T_151,_T_146,_T_136}; // @[HandShaking.scala 741:17]
  assign _T_163 = {out_ready_R_50,out_ready_R_49,out_ready_R_48,out_ready_R_47,out_ready_R_46}; // @[HandShaking.scala 741:17]
  assign _T_169 = {out_ready_R_56,out_ready_R_55,out_ready_R_54,out_ready_R_53,out_ready_R_52,out_ready_R_51,_T_163}; // @[HandShaking.scala 741:17]
  assign _T_174 = {out_ready_R_62,out_ready_R_61,out_ready_R_60,out_ready_R_59,out_ready_R_58,out_ready_R_57}; // @[HandShaking.scala 741:17]
  assign _T_181 = {out_ready_R_68,out_ready_R_67,out_ready_R_66,out_ready_R_65,out_ready_R_64,out_ready_R_63,_T_174,_T_169}; // @[HandShaking.scala 741:17]
  assign _T_186 = {out_ready_R_74,out_ready_R_73,out_ready_R_72,out_ready_R_71,out_ready_R_70,out_ready_R_69}; // @[HandShaking.scala 741:17]
  assign _T_192 = {out_ready_R_80,out_ready_R_79,out_ready_R_78,out_ready_R_77,out_ready_R_76,out_ready_R_75,_T_186}; // @[HandShaking.scala 741:17]
  assign _T_197 = {out_ready_R_86,out_ready_R_85,out_ready_R_84,out_ready_R_83,out_ready_R_82,out_ready_R_81}; // @[HandShaking.scala 741:17]
  assign _T_206 = {out_ready_R_92,out_ready_R_91,out_ready_R_90,out_ready_R_89,out_ready_R_88,out_ready_R_87,_T_197,_T_192,_T_181,_T_159}; // @[HandShaking.scala 741:17]
  assign _T_207 = _T_206 == 93'h1fffffffffffffffffffffff; // @[HandShaking.scala 741:24]
  assign _T_210 = $unsigned(reset); // @[BasicBlock.scala 126:19]
  assign _T_211 = _T_210 == 1'h0; // @[BasicBlock.scala 126:19]
  assign io_MaskBB_0_valid = mask_valid_R_0; // @[HandShaking.scala 726:24]
  assign io_MaskBB_0_bits = {predicate_control_R_1,predicate_control_R_0}; // @[BasicBlock.scala 102:23]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 715:21]
  assign io_Out_0_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 715:21]
  assign io_Out_1_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 715:21]
  assign io_Out_2_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 715:21]
  assign io_Out_3_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 715:21]
  assign io_Out_4_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 715:21]
  assign io_Out_5_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 715:21]
  assign io_Out_6_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 715:21]
  assign io_Out_7_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_8_valid = out_valid_R_8; // @[HandShaking.scala 715:21]
  assign io_Out_8_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_9_valid = out_valid_R_9; // @[HandShaking.scala 715:21]
  assign io_Out_9_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_10_valid = out_valid_R_10; // @[HandShaking.scala 715:21]
  assign io_Out_10_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_11_valid = out_valid_R_11; // @[HandShaking.scala 715:21]
  assign io_Out_11_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_12_valid = out_valid_R_12; // @[HandShaking.scala 715:21]
  assign io_Out_12_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_12_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_13_valid = out_valid_R_13; // @[HandShaking.scala 715:21]
  assign io_Out_13_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_13_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_14_valid = out_valid_R_14; // @[HandShaking.scala 715:21]
  assign io_Out_14_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_14_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_15_valid = out_valid_R_15; // @[HandShaking.scala 715:21]
  assign io_Out_15_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_15_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_16_valid = out_valid_R_16; // @[HandShaking.scala 715:21]
  assign io_Out_16_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_16_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_17_valid = out_valid_R_17; // @[HandShaking.scala 715:21]
  assign io_Out_17_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_17_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_18_valid = out_valid_R_18; // @[HandShaking.scala 715:21]
  assign io_Out_18_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_18_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_19_valid = out_valid_R_19; // @[HandShaking.scala 715:21]
  assign io_Out_19_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_19_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_20_valid = out_valid_R_20; // @[HandShaking.scala 715:21]
  assign io_Out_20_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_20_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_21_valid = out_valid_R_21; // @[HandShaking.scala 715:21]
  assign io_Out_21_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_22_valid = out_valid_R_22; // @[HandShaking.scala 715:21]
  assign io_Out_22_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_22_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_23_valid = out_valid_R_23; // @[HandShaking.scala 715:21]
  assign io_Out_23_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_23_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_24_valid = out_valid_R_24; // @[HandShaking.scala 715:21]
  assign io_Out_24_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_24_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_25_valid = out_valid_R_25; // @[HandShaking.scala 715:21]
  assign io_Out_25_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_25_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_26_valid = out_valid_R_26; // @[HandShaking.scala 715:21]
  assign io_Out_26_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_26_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_27_valid = out_valid_R_27; // @[HandShaking.scala 715:21]
  assign io_Out_27_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_27_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_28_valid = out_valid_R_28; // @[HandShaking.scala 715:21]
  assign io_Out_28_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_28_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_29_valid = out_valid_R_29; // @[HandShaking.scala 715:21]
  assign io_Out_29_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_30_valid = out_valid_R_30; // @[HandShaking.scala 715:21]
  assign io_Out_30_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_30_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_31_valid = out_valid_R_31; // @[HandShaking.scala 715:21]
  assign io_Out_31_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_31_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_32_valid = out_valid_R_32; // @[HandShaking.scala 715:21]
  assign io_Out_32_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_32_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_33_valid = out_valid_R_33; // @[HandShaking.scala 715:21]
  assign io_Out_33_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_33_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_34_valid = out_valid_R_34; // @[HandShaking.scala 715:21]
  assign io_Out_34_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_34_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_35_valid = out_valid_R_35; // @[HandShaking.scala 715:21]
  assign io_Out_35_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_35_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_36_valid = out_valid_R_36; // @[HandShaking.scala 715:21]
  assign io_Out_36_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_36_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_37_valid = out_valid_R_37; // @[HandShaking.scala 715:21]
  assign io_Out_37_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_38_valid = out_valid_R_38; // @[HandShaking.scala 715:21]
  assign io_Out_38_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_38_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_39_valid = out_valid_R_39; // @[HandShaking.scala 715:21]
  assign io_Out_39_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_39_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_40_valid = out_valid_R_40; // @[HandShaking.scala 715:21]
  assign io_Out_40_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_40_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_41_valid = out_valid_R_41; // @[HandShaking.scala 715:21]
  assign io_Out_41_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_41_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_42_valid = out_valid_R_42; // @[HandShaking.scala 715:21]
  assign io_Out_42_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_42_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_43_valid = out_valid_R_43; // @[HandShaking.scala 715:21]
  assign io_Out_43_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_43_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_44_valid = out_valid_R_44; // @[HandShaking.scala 715:21]
  assign io_Out_44_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_44_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_45_valid = out_valid_R_45; // @[HandShaking.scala 715:21]
  assign io_Out_45_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_45_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_46_valid = out_valid_R_46; // @[HandShaking.scala 715:21]
  assign io_Out_46_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_47_valid = out_valid_R_47; // @[HandShaking.scala 715:21]
  assign io_Out_47_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_47_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_48_valid = out_valid_R_48; // @[HandShaking.scala 715:21]
  assign io_Out_48_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_48_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_49_valid = out_valid_R_49; // @[HandShaking.scala 715:21]
  assign io_Out_49_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_49_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_50_valid = out_valid_R_50; // @[HandShaking.scala 715:21]
  assign io_Out_50_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_50_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_51_valid = out_valid_R_51; // @[HandShaking.scala 715:21]
  assign io_Out_51_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_51_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_52_valid = out_valid_R_52; // @[HandShaking.scala 715:21]
  assign io_Out_52_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_52_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_53_valid = out_valid_R_53; // @[HandShaking.scala 715:21]
  assign io_Out_53_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_53_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_54_valid = out_valid_R_54; // @[HandShaking.scala 715:21]
  assign io_Out_54_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_55_valid = out_valid_R_55; // @[HandShaking.scala 715:21]
  assign io_Out_55_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_55_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_56_valid = out_valid_R_56; // @[HandShaking.scala 715:21]
  assign io_Out_56_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_56_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_57_valid = out_valid_R_57; // @[HandShaking.scala 715:21]
  assign io_Out_57_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_57_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_58_valid = out_valid_R_58; // @[HandShaking.scala 715:21]
  assign io_Out_58_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_58_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_59_valid = out_valid_R_59; // @[HandShaking.scala 715:21]
  assign io_Out_59_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_59_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_60_valid = out_valid_R_60; // @[HandShaking.scala 715:21]
  assign io_Out_60_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_60_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_61_valid = out_valid_R_61; // @[HandShaking.scala 715:21]
  assign io_Out_61_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_61_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_62_valid = out_valid_R_62; // @[HandShaking.scala 715:21]
  assign io_Out_62_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_63_valid = out_valid_R_63; // @[HandShaking.scala 715:21]
  assign io_Out_63_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_63_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_64_valid = out_valid_R_64; // @[HandShaking.scala 715:21]
  assign io_Out_64_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_64_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_65_valid = out_valid_R_65; // @[HandShaking.scala 715:21]
  assign io_Out_65_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_65_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_66_valid = out_valid_R_66; // @[HandShaking.scala 715:21]
  assign io_Out_66_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_66_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_67_valid = out_valid_R_67; // @[HandShaking.scala 715:21]
  assign io_Out_67_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_67_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_68_valid = out_valid_R_68; // @[HandShaking.scala 715:21]
  assign io_Out_68_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_68_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_69_valid = out_valid_R_69; // @[HandShaking.scala 715:21]
  assign io_Out_69_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_69_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_70_valid = out_valid_R_70; // @[HandShaking.scala 715:21]
  assign io_Out_70_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_71_valid = out_valid_R_71; // @[HandShaking.scala 715:21]
  assign io_Out_71_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_71_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_72_valid = out_valid_R_72; // @[HandShaking.scala 715:21]
  assign io_Out_72_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_72_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_73_valid = out_valid_R_73; // @[HandShaking.scala 715:21]
  assign io_Out_73_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_73_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_74_valid = out_valid_R_74; // @[HandShaking.scala 715:21]
  assign io_Out_74_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_74_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_75_valid = out_valid_R_75; // @[HandShaking.scala 715:21]
  assign io_Out_75_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_75_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_76_valid = out_valid_R_76; // @[HandShaking.scala 715:21]
  assign io_Out_76_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_76_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_77_valid = out_valid_R_77; // @[HandShaking.scala 715:21]
  assign io_Out_77_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_77_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_78_valid = out_valid_R_78; // @[HandShaking.scala 715:21]
  assign io_Out_78_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_79_valid = out_valid_R_79; // @[HandShaking.scala 715:21]
  assign io_Out_79_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_79_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_80_valid = out_valid_R_80; // @[HandShaking.scala 715:21]
  assign io_Out_80_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_80_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_81_valid = out_valid_R_81; // @[HandShaking.scala 715:21]
  assign io_Out_81_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_81_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_82_valid = out_valid_R_82; // @[HandShaking.scala 715:21]
  assign io_Out_82_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_82_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_83_valid = out_valid_R_83; // @[HandShaking.scala 715:21]
  assign io_Out_83_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_83_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_84_valid = out_valid_R_84; // @[HandShaking.scala 715:21]
  assign io_Out_84_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_84_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_85_valid = out_valid_R_85; // @[HandShaking.scala 715:21]
  assign io_Out_85_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_85_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_86_valid = out_valid_R_86; // @[HandShaking.scala 715:21]
  assign io_Out_86_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_87_valid = out_valid_R_87; // @[HandShaking.scala 715:21]
  assign io_Out_87_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_87_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_88_valid = out_valid_R_88; // @[HandShaking.scala 715:21]
  assign io_Out_88_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_88_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_89_valid = out_valid_R_89; // @[HandShaking.scala 715:21]
  assign io_Out_89_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_89_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_90_valid = out_valid_R_90; // @[HandShaking.scala 715:21]
  assign io_Out_90_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_90_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_91_valid = out_valid_R_91; // @[HandShaking.scala 715:21]
  assign io_Out_91_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_91_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_Out_92_valid = out_valid_R_92; // @[HandShaking.scala 715:21]
  assign io_Out_92_bits_taskID = predicate_in_R_0_taskID | predicate_in_R_1_taskID; // @[BasicBlock.scala 97:27]
  assign io_Out_92_bits_control = predicate_in_R_0_control | predicate_in_R_1_control; // @[BasicBlock.scala 96:28]
  assign io_predicateIn_0_ready = ~ predicate_valid_R_0; // @[BasicBlock.scala 86:29]
  assign io_predicateIn_1_ready = ~ predicate_valid_R_1; // @[BasicBlock.scala 86:29]
  assign _GEN_677 = _T_112 == 1'h0; // @[BasicBlock.scala 126:19]
  assign _GEN_678 = _GEN_677 & state; // @[BasicBlock.scala 126:19]
  assign _GEN_679 = _GEN_678 & _T_207; // @[BasicBlock.scala 126:19]
  assign _GEN_680 = _GEN_679 & predicate; // @[BasicBlock.scala 126:19]
  assign _GEN_684 = predicate == 1'h0; // @[BasicBlock.scala 132:19]
  assign _GEN_685 = _GEN_679 & _GEN_684; // @[BasicBlock.scala 132:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_ready_R_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_ready_R_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_ready_R_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_ready_R_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_ready_R_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_ready_R_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  out_ready_R_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_ready_R_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  out_ready_R_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  out_ready_R_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  out_ready_R_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  out_ready_R_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  out_ready_R_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  out_ready_R_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  out_ready_R_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  out_ready_R_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  out_ready_R_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  out_ready_R_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  out_ready_R_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  out_ready_R_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  out_ready_R_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  out_ready_R_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  out_ready_R_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  out_ready_R_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  out_ready_R_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  out_ready_R_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  out_ready_R_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  out_ready_R_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  out_ready_R_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  out_ready_R_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  out_ready_R_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  out_ready_R_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  out_ready_R_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  out_ready_R_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  out_ready_R_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  out_ready_R_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  out_ready_R_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  out_ready_R_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  out_ready_R_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  out_ready_R_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  out_ready_R_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  out_ready_R_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  out_ready_R_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  out_ready_R_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  out_ready_R_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  out_ready_R_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  out_ready_R_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  out_ready_R_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  out_ready_R_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  out_ready_R_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  out_ready_R_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  out_ready_R_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  out_ready_R_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  out_ready_R_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  out_ready_R_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  out_ready_R_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  out_ready_R_64 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  out_ready_R_65 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  out_ready_R_66 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  out_ready_R_67 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  out_ready_R_68 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  out_ready_R_69 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  out_ready_R_70 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  out_ready_R_71 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  out_ready_R_72 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  out_ready_R_73 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  out_ready_R_74 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  out_ready_R_75 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  out_ready_R_76 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  out_ready_R_77 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  out_ready_R_78 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  out_ready_R_79 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  out_ready_R_80 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  out_ready_R_81 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  out_ready_R_82 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  out_ready_R_83 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  out_ready_R_84 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  out_ready_R_85 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  out_ready_R_86 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  out_ready_R_87 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  out_ready_R_88 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  out_ready_R_89 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  out_ready_R_90 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  out_ready_R_91 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  out_ready_R_92 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  out_valid_R_8 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  out_valid_R_9 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  out_valid_R_10 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  out_valid_R_11 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  out_valid_R_12 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  out_valid_R_13 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  out_valid_R_14 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  out_valid_R_15 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  out_valid_R_16 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  out_valid_R_17 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  out_valid_R_18 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  out_valid_R_19 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  out_valid_R_20 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  out_valid_R_21 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  out_valid_R_22 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  out_valid_R_23 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  out_valid_R_24 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  out_valid_R_25 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  out_valid_R_26 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  out_valid_R_27 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  out_valid_R_28 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  out_valid_R_29 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  out_valid_R_30 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  out_valid_R_31 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  out_valid_R_32 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  out_valid_R_33 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  out_valid_R_34 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  out_valid_R_35 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  out_valid_R_36 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  out_valid_R_37 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  out_valid_R_38 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  out_valid_R_39 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  out_valid_R_40 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  out_valid_R_41 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  out_valid_R_42 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  out_valid_R_43 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  out_valid_R_44 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  out_valid_R_45 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  out_valid_R_46 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  out_valid_R_47 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  out_valid_R_48 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  out_valid_R_49 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  out_valid_R_50 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  out_valid_R_51 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  out_valid_R_52 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  out_valid_R_53 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  out_valid_R_54 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  out_valid_R_55 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  out_valid_R_56 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  out_valid_R_57 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  out_valid_R_58 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  out_valid_R_59 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  out_valid_R_60 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  out_valid_R_61 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  out_valid_R_62 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  out_valid_R_63 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  out_valid_R_64 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  out_valid_R_65 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  out_valid_R_66 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  out_valid_R_67 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  out_valid_R_68 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  out_valid_R_69 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  out_valid_R_70 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  out_valid_R_71 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  out_valid_R_72 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  out_valid_R_73 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  out_valid_R_74 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  out_valid_R_75 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  out_valid_R_76 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  out_valid_R_77 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  out_valid_R_78 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  out_valid_R_79 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  out_valid_R_80 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  out_valid_R_81 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  out_valid_R_82 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  out_valid_R_83 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  out_valid_R_84 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  out_valid_R_85 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  out_valid_R_86 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  out_valid_R_87 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  out_valid_R_88 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  out_valid_R_89 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  out_valid_R_90 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  out_valid_R_91 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  out_valid_R_92 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  mask_valid_R_0 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  value = _RAND_187[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  predicate_in_R_0_taskID = _RAND_188[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  predicate_in_R_0_control = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  predicate_in_R_1_taskID = _RAND_190[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  predicate_in_R_1_control = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  predicate_control_R_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  predicate_control_R_1 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  predicate_valid_R_0 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  predicate_valid_R_1 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  state = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_2) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_3) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_4) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_5) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_6) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_6) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_6) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_7) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_7) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_7) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_8) begin
          out_ready_R_6 <= io_Out_6_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_6 <= 1'h0;
          end else begin
            if (_T_8) begin
              out_ready_R_6 <= io_Out_6_ready;
            end
          end
        end else begin
          if (_T_8) begin
            out_ready_R_6 <= io_Out_6_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_9) begin
          out_ready_R_7 <= io_Out_7_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_7 <= 1'h0;
          end else begin
            if (_T_9) begin
              out_ready_R_7 <= io_Out_7_ready;
            end
          end
        end else begin
          if (_T_9) begin
            out_ready_R_7 <= io_Out_7_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_8 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_10) begin
          out_ready_R_8 <= io_Out_8_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_8 <= 1'h0;
          end else begin
            if (_T_10) begin
              out_ready_R_8 <= io_Out_8_ready;
            end
          end
        end else begin
          if (_T_10) begin
            out_ready_R_8 <= io_Out_8_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_9 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_11) begin
          out_ready_R_9 <= io_Out_9_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_9 <= 1'h0;
          end else begin
            if (_T_11) begin
              out_ready_R_9 <= io_Out_9_ready;
            end
          end
        end else begin
          if (_T_11) begin
            out_ready_R_9 <= io_Out_9_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_10 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_12) begin
          out_ready_R_10 <= io_Out_10_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_10 <= 1'h0;
          end else begin
            if (_T_12) begin
              out_ready_R_10 <= io_Out_10_ready;
            end
          end
        end else begin
          if (_T_12) begin
            out_ready_R_10 <= io_Out_10_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_11 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_13) begin
          out_ready_R_11 <= io_Out_11_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_11 <= 1'h0;
          end else begin
            if (_T_13) begin
              out_ready_R_11 <= io_Out_11_ready;
            end
          end
        end else begin
          if (_T_13) begin
            out_ready_R_11 <= io_Out_11_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_12 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_14) begin
          out_ready_R_12 <= io_Out_12_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_12 <= 1'h0;
          end else begin
            if (_T_14) begin
              out_ready_R_12 <= io_Out_12_ready;
            end
          end
        end else begin
          if (_T_14) begin
            out_ready_R_12 <= io_Out_12_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_13 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_15) begin
          out_ready_R_13 <= io_Out_13_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_13 <= 1'h0;
          end else begin
            if (_T_15) begin
              out_ready_R_13 <= io_Out_13_ready;
            end
          end
        end else begin
          if (_T_15) begin
            out_ready_R_13 <= io_Out_13_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_14 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_16) begin
          out_ready_R_14 <= io_Out_14_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_14 <= 1'h0;
          end else begin
            if (_T_16) begin
              out_ready_R_14 <= io_Out_14_ready;
            end
          end
        end else begin
          if (_T_16) begin
            out_ready_R_14 <= io_Out_14_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_15 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_17) begin
          out_ready_R_15 <= io_Out_15_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_15 <= 1'h0;
          end else begin
            if (_T_17) begin
              out_ready_R_15 <= io_Out_15_ready;
            end
          end
        end else begin
          if (_T_17) begin
            out_ready_R_15 <= io_Out_15_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_16 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_18) begin
          out_ready_R_16 <= io_Out_16_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_16 <= 1'h0;
          end else begin
            if (_T_18) begin
              out_ready_R_16 <= io_Out_16_ready;
            end
          end
        end else begin
          if (_T_18) begin
            out_ready_R_16 <= io_Out_16_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_17 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_19) begin
          out_ready_R_17 <= io_Out_17_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_17 <= 1'h0;
          end else begin
            if (_T_19) begin
              out_ready_R_17 <= io_Out_17_ready;
            end
          end
        end else begin
          if (_T_19) begin
            out_ready_R_17 <= io_Out_17_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_18 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_20) begin
          out_ready_R_18 <= io_Out_18_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_18 <= 1'h0;
          end else begin
            if (_T_20) begin
              out_ready_R_18 <= io_Out_18_ready;
            end
          end
        end else begin
          if (_T_20) begin
            out_ready_R_18 <= io_Out_18_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_19 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_21) begin
          out_ready_R_19 <= io_Out_19_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_19 <= 1'h0;
          end else begin
            if (_T_21) begin
              out_ready_R_19 <= io_Out_19_ready;
            end
          end
        end else begin
          if (_T_21) begin
            out_ready_R_19 <= io_Out_19_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_20 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_22) begin
          out_ready_R_20 <= io_Out_20_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_20 <= 1'h0;
          end else begin
            if (_T_22) begin
              out_ready_R_20 <= io_Out_20_ready;
            end
          end
        end else begin
          if (_T_22) begin
            out_ready_R_20 <= io_Out_20_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_21 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_23) begin
          out_ready_R_21 <= io_Out_21_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_21 <= 1'h0;
          end else begin
            if (_T_23) begin
              out_ready_R_21 <= io_Out_21_ready;
            end
          end
        end else begin
          if (_T_23) begin
            out_ready_R_21 <= io_Out_21_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_22 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_24) begin
          out_ready_R_22 <= io_Out_22_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_22 <= 1'h0;
          end else begin
            if (_T_24) begin
              out_ready_R_22 <= io_Out_22_ready;
            end
          end
        end else begin
          if (_T_24) begin
            out_ready_R_22 <= io_Out_22_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_23 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_25) begin
          out_ready_R_23 <= io_Out_23_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_23 <= 1'h0;
          end else begin
            if (_T_25) begin
              out_ready_R_23 <= io_Out_23_ready;
            end
          end
        end else begin
          if (_T_25) begin
            out_ready_R_23 <= io_Out_23_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_24 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_26) begin
          out_ready_R_24 <= io_Out_24_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_24 <= 1'h0;
          end else begin
            if (_T_26) begin
              out_ready_R_24 <= io_Out_24_ready;
            end
          end
        end else begin
          if (_T_26) begin
            out_ready_R_24 <= io_Out_24_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_25 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_27) begin
          out_ready_R_25 <= io_Out_25_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_25 <= 1'h0;
          end else begin
            if (_T_27) begin
              out_ready_R_25 <= io_Out_25_ready;
            end
          end
        end else begin
          if (_T_27) begin
            out_ready_R_25 <= io_Out_25_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_26 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_28) begin
          out_ready_R_26 <= io_Out_26_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_26 <= 1'h0;
          end else begin
            if (_T_28) begin
              out_ready_R_26 <= io_Out_26_ready;
            end
          end
        end else begin
          if (_T_28) begin
            out_ready_R_26 <= io_Out_26_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_27 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_29) begin
          out_ready_R_27 <= io_Out_27_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_27 <= 1'h0;
          end else begin
            if (_T_29) begin
              out_ready_R_27 <= io_Out_27_ready;
            end
          end
        end else begin
          if (_T_29) begin
            out_ready_R_27 <= io_Out_27_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_28 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_30) begin
          out_ready_R_28 <= io_Out_28_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_28 <= 1'h0;
          end else begin
            if (_T_30) begin
              out_ready_R_28 <= io_Out_28_ready;
            end
          end
        end else begin
          if (_T_30) begin
            out_ready_R_28 <= io_Out_28_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_29 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_31) begin
          out_ready_R_29 <= io_Out_29_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_29 <= 1'h0;
          end else begin
            if (_T_31) begin
              out_ready_R_29 <= io_Out_29_ready;
            end
          end
        end else begin
          if (_T_31) begin
            out_ready_R_29 <= io_Out_29_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_30 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_32) begin
          out_ready_R_30 <= io_Out_30_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_30 <= 1'h0;
          end else begin
            if (_T_32) begin
              out_ready_R_30 <= io_Out_30_ready;
            end
          end
        end else begin
          if (_T_32) begin
            out_ready_R_30 <= io_Out_30_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_31 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_33) begin
          out_ready_R_31 <= io_Out_31_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_31 <= 1'h0;
          end else begin
            if (_T_33) begin
              out_ready_R_31 <= io_Out_31_ready;
            end
          end
        end else begin
          if (_T_33) begin
            out_ready_R_31 <= io_Out_31_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_32 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_34) begin
          out_ready_R_32 <= io_Out_32_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_32 <= 1'h0;
          end else begin
            if (_T_34) begin
              out_ready_R_32 <= io_Out_32_ready;
            end
          end
        end else begin
          if (_T_34) begin
            out_ready_R_32 <= io_Out_32_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_33 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_35) begin
          out_ready_R_33 <= io_Out_33_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_33 <= 1'h0;
          end else begin
            if (_T_35) begin
              out_ready_R_33 <= io_Out_33_ready;
            end
          end
        end else begin
          if (_T_35) begin
            out_ready_R_33 <= io_Out_33_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_34 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_36) begin
          out_ready_R_34 <= io_Out_34_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_34 <= 1'h0;
          end else begin
            if (_T_36) begin
              out_ready_R_34 <= io_Out_34_ready;
            end
          end
        end else begin
          if (_T_36) begin
            out_ready_R_34 <= io_Out_34_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_35 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_37) begin
          out_ready_R_35 <= io_Out_35_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_35 <= 1'h0;
          end else begin
            if (_T_37) begin
              out_ready_R_35 <= io_Out_35_ready;
            end
          end
        end else begin
          if (_T_37) begin
            out_ready_R_35 <= io_Out_35_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_36 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_38) begin
          out_ready_R_36 <= io_Out_36_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_36 <= 1'h0;
          end else begin
            if (_T_38) begin
              out_ready_R_36 <= io_Out_36_ready;
            end
          end
        end else begin
          if (_T_38) begin
            out_ready_R_36 <= io_Out_36_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_37 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_39) begin
          out_ready_R_37 <= io_Out_37_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_37 <= 1'h0;
          end else begin
            if (_T_39) begin
              out_ready_R_37 <= io_Out_37_ready;
            end
          end
        end else begin
          if (_T_39) begin
            out_ready_R_37 <= io_Out_37_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_38 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_40) begin
          out_ready_R_38 <= io_Out_38_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_38 <= 1'h0;
          end else begin
            if (_T_40) begin
              out_ready_R_38 <= io_Out_38_ready;
            end
          end
        end else begin
          if (_T_40) begin
            out_ready_R_38 <= io_Out_38_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_39 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_41) begin
          out_ready_R_39 <= io_Out_39_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_39 <= 1'h0;
          end else begin
            if (_T_41) begin
              out_ready_R_39 <= io_Out_39_ready;
            end
          end
        end else begin
          if (_T_41) begin
            out_ready_R_39 <= io_Out_39_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_40 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_42) begin
          out_ready_R_40 <= io_Out_40_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_40 <= 1'h0;
          end else begin
            if (_T_42) begin
              out_ready_R_40 <= io_Out_40_ready;
            end
          end
        end else begin
          if (_T_42) begin
            out_ready_R_40 <= io_Out_40_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_41 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_43) begin
          out_ready_R_41 <= io_Out_41_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_41 <= 1'h0;
          end else begin
            if (_T_43) begin
              out_ready_R_41 <= io_Out_41_ready;
            end
          end
        end else begin
          if (_T_43) begin
            out_ready_R_41 <= io_Out_41_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_42 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_44) begin
          out_ready_R_42 <= io_Out_42_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_42 <= 1'h0;
          end else begin
            if (_T_44) begin
              out_ready_R_42 <= io_Out_42_ready;
            end
          end
        end else begin
          if (_T_44) begin
            out_ready_R_42 <= io_Out_42_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_43 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_45) begin
          out_ready_R_43 <= io_Out_43_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_43 <= 1'h0;
          end else begin
            if (_T_45) begin
              out_ready_R_43 <= io_Out_43_ready;
            end
          end
        end else begin
          if (_T_45) begin
            out_ready_R_43 <= io_Out_43_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_44 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_46) begin
          out_ready_R_44 <= io_Out_44_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_44 <= 1'h0;
          end else begin
            if (_T_46) begin
              out_ready_R_44 <= io_Out_44_ready;
            end
          end
        end else begin
          if (_T_46) begin
            out_ready_R_44 <= io_Out_44_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_45 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_47) begin
          out_ready_R_45 <= io_Out_45_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_45 <= 1'h0;
          end else begin
            if (_T_47) begin
              out_ready_R_45 <= io_Out_45_ready;
            end
          end
        end else begin
          if (_T_47) begin
            out_ready_R_45 <= io_Out_45_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_46 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_48) begin
          out_ready_R_46 <= io_Out_46_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_46 <= 1'h0;
          end else begin
            if (_T_48) begin
              out_ready_R_46 <= io_Out_46_ready;
            end
          end
        end else begin
          if (_T_48) begin
            out_ready_R_46 <= io_Out_46_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_47 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_49) begin
          out_ready_R_47 <= io_Out_47_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_47 <= 1'h0;
          end else begin
            if (_T_49) begin
              out_ready_R_47 <= io_Out_47_ready;
            end
          end
        end else begin
          if (_T_49) begin
            out_ready_R_47 <= io_Out_47_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_48 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_50) begin
          out_ready_R_48 <= io_Out_48_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_48 <= 1'h0;
          end else begin
            if (_T_50) begin
              out_ready_R_48 <= io_Out_48_ready;
            end
          end
        end else begin
          if (_T_50) begin
            out_ready_R_48 <= io_Out_48_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_49 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_51) begin
          out_ready_R_49 <= io_Out_49_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_49 <= 1'h0;
          end else begin
            if (_T_51) begin
              out_ready_R_49 <= io_Out_49_ready;
            end
          end
        end else begin
          if (_T_51) begin
            out_ready_R_49 <= io_Out_49_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_50 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_52) begin
          out_ready_R_50 <= io_Out_50_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_50 <= 1'h0;
          end else begin
            if (_T_52) begin
              out_ready_R_50 <= io_Out_50_ready;
            end
          end
        end else begin
          if (_T_52) begin
            out_ready_R_50 <= io_Out_50_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_51 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_53) begin
          out_ready_R_51 <= io_Out_51_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_51 <= 1'h0;
          end else begin
            if (_T_53) begin
              out_ready_R_51 <= io_Out_51_ready;
            end
          end
        end else begin
          if (_T_53) begin
            out_ready_R_51 <= io_Out_51_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_52 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_54) begin
          out_ready_R_52 <= io_Out_52_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_52 <= 1'h0;
          end else begin
            if (_T_54) begin
              out_ready_R_52 <= io_Out_52_ready;
            end
          end
        end else begin
          if (_T_54) begin
            out_ready_R_52 <= io_Out_52_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_53 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_55) begin
          out_ready_R_53 <= io_Out_53_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_53 <= 1'h0;
          end else begin
            if (_T_55) begin
              out_ready_R_53 <= io_Out_53_ready;
            end
          end
        end else begin
          if (_T_55) begin
            out_ready_R_53 <= io_Out_53_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_54 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_56) begin
          out_ready_R_54 <= io_Out_54_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_54 <= 1'h0;
          end else begin
            if (_T_56) begin
              out_ready_R_54 <= io_Out_54_ready;
            end
          end
        end else begin
          if (_T_56) begin
            out_ready_R_54 <= io_Out_54_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_55 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_57) begin
          out_ready_R_55 <= io_Out_55_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_55 <= 1'h0;
          end else begin
            if (_T_57) begin
              out_ready_R_55 <= io_Out_55_ready;
            end
          end
        end else begin
          if (_T_57) begin
            out_ready_R_55 <= io_Out_55_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_56 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_58) begin
          out_ready_R_56 <= io_Out_56_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_56 <= 1'h0;
          end else begin
            if (_T_58) begin
              out_ready_R_56 <= io_Out_56_ready;
            end
          end
        end else begin
          if (_T_58) begin
            out_ready_R_56 <= io_Out_56_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_57 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_59) begin
          out_ready_R_57 <= io_Out_57_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_57 <= 1'h0;
          end else begin
            if (_T_59) begin
              out_ready_R_57 <= io_Out_57_ready;
            end
          end
        end else begin
          if (_T_59) begin
            out_ready_R_57 <= io_Out_57_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_58 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_60) begin
          out_ready_R_58 <= io_Out_58_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_58 <= 1'h0;
          end else begin
            if (_T_60) begin
              out_ready_R_58 <= io_Out_58_ready;
            end
          end
        end else begin
          if (_T_60) begin
            out_ready_R_58 <= io_Out_58_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_59 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_61) begin
          out_ready_R_59 <= io_Out_59_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_59 <= 1'h0;
          end else begin
            if (_T_61) begin
              out_ready_R_59 <= io_Out_59_ready;
            end
          end
        end else begin
          if (_T_61) begin
            out_ready_R_59 <= io_Out_59_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_60 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_62) begin
          out_ready_R_60 <= io_Out_60_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_60 <= 1'h0;
          end else begin
            if (_T_62) begin
              out_ready_R_60 <= io_Out_60_ready;
            end
          end
        end else begin
          if (_T_62) begin
            out_ready_R_60 <= io_Out_60_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_61 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_63) begin
          out_ready_R_61 <= io_Out_61_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_61 <= 1'h0;
          end else begin
            if (_T_63) begin
              out_ready_R_61 <= io_Out_61_ready;
            end
          end
        end else begin
          if (_T_63) begin
            out_ready_R_61 <= io_Out_61_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_62 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_64) begin
          out_ready_R_62 <= io_Out_62_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_62 <= 1'h0;
          end else begin
            if (_T_64) begin
              out_ready_R_62 <= io_Out_62_ready;
            end
          end
        end else begin
          if (_T_64) begin
            out_ready_R_62 <= io_Out_62_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_63 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_65) begin
          out_ready_R_63 <= io_Out_63_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_63 <= 1'h0;
          end else begin
            if (_T_65) begin
              out_ready_R_63 <= io_Out_63_ready;
            end
          end
        end else begin
          if (_T_65) begin
            out_ready_R_63 <= io_Out_63_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_64 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_66) begin
          out_ready_R_64 <= io_Out_64_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_64 <= 1'h0;
          end else begin
            if (_T_66) begin
              out_ready_R_64 <= io_Out_64_ready;
            end
          end
        end else begin
          if (_T_66) begin
            out_ready_R_64 <= io_Out_64_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_65 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_67) begin
          out_ready_R_65 <= io_Out_65_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_65 <= 1'h0;
          end else begin
            if (_T_67) begin
              out_ready_R_65 <= io_Out_65_ready;
            end
          end
        end else begin
          if (_T_67) begin
            out_ready_R_65 <= io_Out_65_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_66 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_68) begin
          out_ready_R_66 <= io_Out_66_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_66 <= 1'h0;
          end else begin
            if (_T_68) begin
              out_ready_R_66 <= io_Out_66_ready;
            end
          end
        end else begin
          if (_T_68) begin
            out_ready_R_66 <= io_Out_66_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_67 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_69) begin
          out_ready_R_67 <= io_Out_67_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_67 <= 1'h0;
          end else begin
            if (_T_69) begin
              out_ready_R_67 <= io_Out_67_ready;
            end
          end
        end else begin
          if (_T_69) begin
            out_ready_R_67 <= io_Out_67_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_68 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_70) begin
          out_ready_R_68 <= io_Out_68_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_68 <= 1'h0;
          end else begin
            if (_T_70) begin
              out_ready_R_68 <= io_Out_68_ready;
            end
          end
        end else begin
          if (_T_70) begin
            out_ready_R_68 <= io_Out_68_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_69 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_71) begin
          out_ready_R_69 <= io_Out_69_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_69 <= 1'h0;
          end else begin
            if (_T_71) begin
              out_ready_R_69 <= io_Out_69_ready;
            end
          end
        end else begin
          if (_T_71) begin
            out_ready_R_69 <= io_Out_69_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_70 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_72) begin
          out_ready_R_70 <= io_Out_70_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_70 <= 1'h0;
          end else begin
            if (_T_72) begin
              out_ready_R_70 <= io_Out_70_ready;
            end
          end
        end else begin
          if (_T_72) begin
            out_ready_R_70 <= io_Out_70_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_71 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_73) begin
          out_ready_R_71 <= io_Out_71_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_71 <= 1'h0;
          end else begin
            if (_T_73) begin
              out_ready_R_71 <= io_Out_71_ready;
            end
          end
        end else begin
          if (_T_73) begin
            out_ready_R_71 <= io_Out_71_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_72 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_74) begin
          out_ready_R_72 <= io_Out_72_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_72 <= 1'h0;
          end else begin
            if (_T_74) begin
              out_ready_R_72 <= io_Out_72_ready;
            end
          end
        end else begin
          if (_T_74) begin
            out_ready_R_72 <= io_Out_72_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_73 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_75) begin
          out_ready_R_73 <= io_Out_73_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_73 <= 1'h0;
          end else begin
            if (_T_75) begin
              out_ready_R_73 <= io_Out_73_ready;
            end
          end
        end else begin
          if (_T_75) begin
            out_ready_R_73 <= io_Out_73_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_74 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_76) begin
          out_ready_R_74 <= io_Out_74_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_74 <= 1'h0;
          end else begin
            if (_T_76) begin
              out_ready_R_74 <= io_Out_74_ready;
            end
          end
        end else begin
          if (_T_76) begin
            out_ready_R_74 <= io_Out_74_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_75 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_77) begin
          out_ready_R_75 <= io_Out_75_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_75 <= 1'h0;
          end else begin
            if (_T_77) begin
              out_ready_R_75 <= io_Out_75_ready;
            end
          end
        end else begin
          if (_T_77) begin
            out_ready_R_75 <= io_Out_75_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_76 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_78) begin
          out_ready_R_76 <= io_Out_76_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_76 <= 1'h0;
          end else begin
            if (_T_78) begin
              out_ready_R_76 <= io_Out_76_ready;
            end
          end
        end else begin
          if (_T_78) begin
            out_ready_R_76 <= io_Out_76_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_77 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_79) begin
          out_ready_R_77 <= io_Out_77_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_77 <= 1'h0;
          end else begin
            if (_T_79) begin
              out_ready_R_77 <= io_Out_77_ready;
            end
          end
        end else begin
          if (_T_79) begin
            out_ready_R_77 <= io_Out_77_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_78 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_80) begin
          out_ready_R_78 <= io_Out_78_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_78 <= 1'h0;
          end else begin
            if (_T_80) begin
              out_ready_R_78 <= io_Out_78_ready;
            end
          end
        end else begin
          if (_T_80) begin
            out_ready_R_78 <= io_Out_78_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_79 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_81) begin
          out_ready_R_79 <= io_Out_79_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_79 <= 1'h0;
          end else begin
            if (_T_81) begin
              out_ready_R_79 <= io_Out_79_ready;
            end
          end
        end else begin
          if (_T_81) begin
            out_ready_R_79 <= io_Out_79_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_80 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_82) begin
          out_ready_R_80 <= io_Out_80_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_80 <= 1'h0;
          end else begin
            if (_T_82) begin
              out_ready_R_80 <= io_Out_80_ready;
            end
          end
        end else begin
          if (_T_82) begin
            out_ready_R_80 <= io_Out_80_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_81 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_83) begin
          out_ready_R_81 <= io_Out_81_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_81 <= 1'h0;
          end else begin
            if (_T_83) begin
              out_ready_R_81 <= io_Out_81_ready;
            end
          end
        end else begin
          if (_T_83) begin
            out_ready_R_81 <= io_Out_81_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_82 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_84) begin
          out_ready_R_82 <= io_Out_82_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_82 <= 1'h0;
          end else begin
            if (_T_84) begin
              out_ready_R_82 <= io_Out_82_ready;
            end
          end
        end else begin
          if (_T_84) begin
            out_ready_R_82 <= io_Out_82_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_83 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_85) begin
          out_ready_R_83 <= io_Out_83_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_83 <= 1'h0;
          end else begin
            if (_T_85) begin
              out_ready_R_83 <= io_Out_83_ready;
            end
          end
        end else begin
          if (_T_85) begin
            out_ready_R_83 <= io_Out_83_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_84 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_86) begin
          out_ready_R_84 <= io_Out_84_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_84 <= 1'h0;
          end else begin
            if (_T_86) begin
              out_ready_R_84 <= io_Out_84_ready;
            end
          end
        end else begin
          if (_T_86) begin
            out_ready_R_84 <= io_Out_84_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_85 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_87) begin
          out_ready_R_85 <= io_Out_85_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_85 <= 1'h0;
          end else begin
            if (_T_87) begin
              out_ready_R_85 <= io_Out_85_ready;
            end
          end
        end else begin
          if (_T_87) begin
            out_ready_R_85 <= io_Out_85_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_86 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_88) begin
          out_ready_R_86 <= io_Out_86_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_86 <= 1'h0;
          end else begin
            if (_T_88) begin
              out_ready_R_86 <= io_Out_86_ready;
            end
          end
        end else begin
          if (_T_88) begin
            out_ready_R_86 <= io_Out_86_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_87 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_89) begin
          out_ready_R_87 <= io_Out_87_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_87 <= 1'h0;
          end else begin
            if (_T_89) begin
              out_ready_R_87 <= io_Out_87_ready;
            end
          end
        end else begin
          if (_T_89) begin
            out_ready_R_87 <= io_Out_87_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_88 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_90) begin
          out_ready_R_88 <= io_Out_88_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_88 <= 1'h0;
          end else begin
            if (_T_90) begin
              out_ready_R_88 <= io_Out_88_ready;
            end
          end
        end else begin
          if (_T_90) begin
            out_ready_R_88 <= io_Out_88_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_89 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_91) begin
          out_ready_R_89 <= io_Out_89_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_89 <= 1'h0;
          end else begin
            if (_T_91) begin
              out_ready_R_89 <= io_Out_89_ready;
            end
          end
        end else begin
          if (_T_91) begin
            out_ready_R_89 <= io_Out_89_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_90 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_92) begin
          out_ready_R_90 <= io_Out_90_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_90 <= 1'h0;
          end else begin
            if (_T_92) begin
              out_ready_R_90 <= io_Out_90_ready;
            end
          end
        end else begin
          if (_T_92) begin
            out_ready_R_90 <= io_Out_90_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_91 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_93) begin
          out_ready_R_91 <= io_Out_91_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_91 <= 1'h0;
          end else begin
            if (_T_93) begin
              out_ready_R_91 <= io_Out_91_ready;
            end
          end
        end else begin
          if (_T_93) begin
            out_ready_R_91 <= io_Out_91_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_92 <= 1'h0;
    end else begin
      if (_T_112) begin
        if (_T_94) begin
          out_ready_R_92 <= io_Out_92_ready;
        end
      end else begin
        if (state) begin
          if (_T_207) begin
            out_ready_R_92 <= 1'h0;
          end else begin
            if (_T_94) begin
              out_ready_R_92 <= io_Out_92_ready;
            end
          end
        end else begin
          if (_T_94) begin
            out_ready_R_92 <= io_Out_92_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_0 <= _GEN_197;
      end else begin
        if (_T_2) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_1 <= _GEN_198;
      end else begin
        if (_T_3) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_2 <= _GEN_199;
      end else begin
        if (_T_4) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_3 <= _GEN_200;
      end else begin
        if (_T_5) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_4 <= _GEN_201;
      end else begin
        if (_T_6) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_5 <= _GEN_202;
      end else begin
        if (_T_7) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_6 <= _GEN_203;
      end else begin
        if (_T_8) begin
          out_valid_R_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_7 <= _GEN_204;
      end else begin
        if (_T_9) begin
          out_valid_R_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_8 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_8 <= _GEN_205;
      end else begin
        if (_T_10) begin
          out_valid_R_8 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_9 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_9 <= _GEN_206;
      end else begin
        if (_T_11) begin
          out_valid_R_9 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_10 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_10 <= _GEN_207;
      end else begin
        if (_T_12) begin
          out_valid_R_10 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_11 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_11 <= _GEN_208;
      end else begin
        if (_T_13) begin
          out_valid_R_11 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_12 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_12 <= _GEN_209;
      end else begin
        if (_T_14) begin
          out_valid_R_12 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_13 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_13 <= _GEN_210;
      end else begin
        if (_T_15) begin
          out_valid_R_13 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_14 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_14 <= _GEN_211;
      end else begin
        if (_T_16) begin
          out_valid_R_14 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_15 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_15 <= _GEN_212;
      end else begin
        if (_T_17) begin
          out_valid_R_15 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_16 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_16 <= _GEN_213;
      end else begin
        if (_T_18) begin
          out_valid_R_16 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_17 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_17 <= _GEN_214;
      end else begin
        if (_T_19) begin
          out_valid_R_17 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_18 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_18 <= _GEN_215;
      end else begin
        if (_T_20) begin
          out_valid_R_18 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_19 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_19 <= _GEN_216;
      end else begin
        if (_T_21) begin
          out_valid_R_19 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_20 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_20 <= _GEN_217;
      end else begin
        if (_T_22) begin
          out_valid_R_20 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_21 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_21 <= _GEN_218;
      end else begin
        if (_T_23) begin
          out_valid_R_21 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_22 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_22 <= _GEN_219;
      end else begin
        if (_T_24) begin
          out_valid_R_22 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_23 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_23 <= _GEN_220;
      end else begin
        if (_T_25) begin
          out_valid_R_23 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_24 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_24 <= _GEN_221;
      end else begin
        if (_T_26) begin
          out_valid_R_24 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_25 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_25 <= _GEN_222;
      end else begin
        if (_T_27) begin
          out_valid_R_25 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_26 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_26 <= _GEN_223;
      end else begin
        if (_T_28) begin
          out_valid_R_26 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_27 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_27 <= _GEN_224;
      end else begin
        if (_T_29) begin
          out_valid_R_27 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_28 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_28 <= _GEN_225;
      end else begin
        if (_T_30) begin
          out_valid_R_28 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_29 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_29 <= _GEN_226;
      end else begin
        if (_T_31) begin
          out_valid_R_29 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_30 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_30 <= _GEN_227;
      end else begin
        if (_T_32) begin
          out_valid_R_30 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_31 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_31 <= _GEN_228;
      end else begin
        if (_T_33) begin
          out_valid_R_31 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_32 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_32 <= _GEN_229;
      end else begin
        if (_T_34) begin
          out_valid_R_32 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_33 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_33 <= _GEN_230;
      end else begin
        if (_T_35) begin
          out_valid_R_33 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_34 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_34 <= _GEN_231;
      end else begin
        if (_T_36) begin
          out_valid_R_34 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_35 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_35 <= _GEN_232;
      end else begin
        if (_T_37) begin
          out_valid_R_35 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_36 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_36 <= _GEN_233;
      end else begin
        if (_T_38) begin
          out_valid_R_36 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_37 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_37 <= _GEN_234;
      end else begin
        if (_T_39) begin
          out_valid_R_37 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_38 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_38 <= _GEN_235;
      end else begin
        if (_T_40) begin
          out_valid_R_38 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_39 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_39 <= _GEN_236;
      end else begin
        if (_T_41) begin
          out_valid_R_39 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_40 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_40 <= _GEN_237;
      end else begin
        if (_T_42) begin
          out_valid_R_40 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_41 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_41 <= _GEN_238;
      end else begin
        if (_T_43) begin
          out_valid_R_41 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_42 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_42 <= _GEN_239;
      end else begin
        if (_T_44) begin
          out_valid_R_42 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_43 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_43 <= _GEN_240;
      end else begin
        if (_T_45) begin
          out_valid_R_43 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_44 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_44 <= _GEN_241;
      end else begin
        if (_T_46) begin
          out_valid_R_44 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_45 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_45 <= _GEN_242;
      end else begin
        if (_T_47) begin
          out_valid_R_45 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_46 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_46 <= _GEN_243;
      end else begin
        if (_T_48) begin
          out_valid_R_46 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_47 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_47 <= _GEN_244;
      end else begin
        if (_T_49) begin
          out_valid_R_47 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_48 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_48 <= _GEN_245;
      end else begin
        if (_T_50) begin
          out_valid_R_48 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_49 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_49 <= _GEN_246;
      end else begin
        if (_T_51) begin
          out_valid_R_49 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_50 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_50 <= _GEN_247;
      end else begin
        if (_T_52) begin
          out_valid_R_50 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_51 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_51 <= _GEN_248;
      end else begin
        if (_T_53) begin
          out_valid_R_51 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_52 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_52 <= _GEN_249;
      end else begin
        if (_T_54) begin
          out_valid_R_52 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_53 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_53 <= _GEN_250;
      end else begin
        if (_T_55) begin
          out_valid_R_53 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_54 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_54 <= _GEN_251;
      end else begin
        if (_T_56) begin
          out_valid_R_54 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_55 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_55 <= _GEN_252;
      end else begin
        if (_T_57) begin
          out_valid_R_55 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_56 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_56 <= _GEN_253;
      end else begin
        if (_T_58) begin
          out_valid_R_56 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_57 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_57 <= _GEN_254;
      end else begin
        if (_T_59) begin
          out_valid_R_57 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_58 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_58 <= _GEN_255;
      end else begin
        if (_T_60) begin
          out_valid_R_58 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_59 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_59 <= _GEN_256;
      end else begin
        if (_T_61) begin
          out_valid_R_59 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_60 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_60 <= _GEN_257;
      end else begin
        if (_T_62) begin
          out_valid_R_60 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_61 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_61 <= _GEN_258;
      end else begin
        if (_T_63) begin
          out_valid_R_61 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_62 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_62 <= _GEN_259;
      end else begin
        if (_T_64) begin
          out_valid_R_62 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_63 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_63 <= _GEN_260;
      end else begin
        if (_T_65) begin
          out_valid_R_63 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_64 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_64 <= _GEN_261;
      end else begin
        if (_T_66) begin
          out_valid_R_64 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_65 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_65 <= _GEN_262;
      end else begin
        if (_T_67) begin
          out_valid_R_65 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_66 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_66 <= _GEN_263;
      end else begin
        if (_T_68) begin
          out_valid_R_66 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_67 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_67 <= _GEN_264;
      end else begin
        if (_T_69) begin
          out_valid_R_67 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_68 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_68 <= _GEN_265;
      end else begin
        if (_T_70) begin
          out_valid_R_68 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_69 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_69 <= _GEN_266;
      end else begin
        if (_T_71) begin
          out_valid_R_69 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_70 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_70 <= _GEN_267;
      end else begin
        if (_T_72) begin
          out_valid_R_70 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_71 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_71 <= _GEN_268;
      end else begin
        if (_T_73) begin
          out_valid_R_71 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_72 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_72 <= _GEN_269;
      end else begin
        if (_T_74) begin
          out_valid_R_72 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_73 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_73 <= _GEN_270;
      end else begin
        if (_T_75) begin
          out_valid_R_73 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_74 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_74 <= _GEN_271;
      end else begin
        if (_T_76) begin
          out_valid_R_74 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_75 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_75 <= _GEN_272;
      end else begin
        if (_T_77) begin
          out_valid_R_75 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_76 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_76 <= _GEN_273;
      end else begin
        if (_T_78) begin
          out_valid_R_76 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_77 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_77 <= _GEN_274;
      end else begin
        if (_T_79) begin
          out_valid_R_77 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_78 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_78 <= _GEN_275;
      end else begin
        if (_T_80) begin
          out_valid_R_78 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_79 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_79 <= _GEN_276;
      end else begin
        if (_T_81) begin
          out_valid_R_79 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_80 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_80 <= _GEN_277;
      end else begin
        if (_T_82) begin
          out_valid_R_80 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_81 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_81 <= _GEN_278;
      end else begin
        if (_T_83) begin
          out_valid_R_81 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_82 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_82 <= _GEN_279;
      end else begin
        if (_T_84) begin
          out_valid_R_82 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_83 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_83 <= _GEN_280;
      end else begin
        if (_T_85) begin
          out_valid_R_83 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_84 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_84 <= _GEN_281;
      end else begin
        if (_T_86) begin
          out_valid_R_84 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_85 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_85 <= _GEN_282;
      end else begin
        if (_T_87) begin
          out_valid_R_85 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_86 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_86 <= _GEN_283;
      end else begin
        if (_T_88) begin
          out_valid_R_86 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_87 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_87 <= _GEN_284;
      end else begin
        if (_T_89) begin
          out_valid_R_87 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_88 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_88 <= _GEN_285;
      end else begin
        if (_T_90) begin
          out_valid_R_88 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_89 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_89 <= _GEN_286;
      end else begin
        if (_T_91) begin
          out_valid_R_89 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_90 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_90 <= _GEN_287;
      end else begin
        if (_T_92) begin
          out_valid_R_90 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_91 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_91 <= _GEN_288;
      end else begin
        if (_T_93) begin
          out_valid_R_91 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_92 <= 1'h0;
    end else begin
      if (_T_112) begin
        out_valid_R_92 <= _GEN_289;
      end else begin
        if (_T_94) begin
          out_valid_R_92 <= 1'h0;
        end
      end
    end
    if (reset) begin
      mask_valid_R_0 <= 1'h0;
    end else begin
      if (_T_112) begin
        mask_valid_R_0 <= _GEN_290;
      end else begin
        if (_T_95) begin
          mask_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_98;
    end
    if (reset) begin
      predicate_in_R_0_taskID <= 5'h0;
    end else begin
      if (_T_103) begin
        predicate_in_R_0_taskID <= io_predicateIn_0_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_0_control <= 1'h0;
    end else begin
      if (_T_103) begin
        predicate_in_R_0_control <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_in_R_1_taskID <= 5'h0;
    end else begin
      if (_T_104) begin
        predicate_in_R_1_taskID <= io_predicateIn_1_bits_taskID;
      end
    end
    if (reset) begin
      predicate_in_R_1_control <= 1'h0;
    end else begin
      if (_T_104) begin
        predicate_in_R_1_control <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_0 <= 1'h0;
    end else begin
      if (_T_103) begin
        predicate_control_R_0 <= io_predicateIn_0_bits_control;
      end
    end
    if (reset) begin
      predicate_control_R_1 <= 1'h0;
    end else begin
      if (_T_104) begin
        predicate_control_R_1 <= io_predicateIn_1_bits_control;
      end
    end
    if (reset) begin
      predicate_valid_R_0 <= 1'h0;
    end else begin
      if (_T_112) begin
        predicate_valid_R_0 <= _T_105;
      end else begin
        if (state) begin
          if (_T_207) begin
            predicate_valid_R_0 <= 1'h0;
          end else begin
            predicate_valid_R_0 <= _T_105;
          end
        end else begin
          predicate_valid_R_0 <= _T_105;
        end
      end
    end
    if (reset) begin
      predicate_valid_R_1 <= 1'h0;
    end else begin
      if (_T_112) begin
        predicate_valid_R_1 <= _T_106;
      end else begin
        if (state) begin
          if (_T_207) begin
            predicate_valid_R_1 <= 1'h0;
          end else begin
            predicate_valid_R_1 <= _T_106;
          end
        end else begin
          predicate_valid_R_1 <= _T_106;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_112) begin
        state <= _GEN_291;
      end else begin
        if (state) begin
          if (_T_207) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_680 & _T_211) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [BB]   bb_for_body124: Output fired @ %d, Mask: %d\n",predicate_task,value,_T_111); // @[BasicBlock.scala 126:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_685 & _T_211) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] bb_for_body124: Output fired @ %d -> 0 predicate\n",value); // @[BasicBlock.scala 132:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire [63:0] _T_24; // @[Alu.scala 195:32]
  assign _T_24 = io_in1 * io_in2; // @[Alu.scala 195:32]
  assign io_out = _T_24[31:0]; // @[Alu.scala 236:10]
endmodule
module ComputeNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul0: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_1(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  assign io_out = io_in1 + io_in2; // @[Alu.scala 236:10]
endmodule
module ComputeNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add1: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= 32'h1;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= 32'h1;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= 32'h1;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx252: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= 32'h2;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= 32'h2;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= 32'h2;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx383: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= 32'h3;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= 32'h3;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= 32'h3;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx514: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= 32'h4;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= 32'h4;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= 32'h4;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx625: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= 32'h5;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= 32'h5;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= 32'h5;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx746: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= 32'h6;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= 32'h6;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= 32'h6;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx867: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_6(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= 32'h7;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= 32'h7;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= 32'h7;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx978: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_7(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= 32'h8;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= 32'h8;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= 32'h8;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx1099: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [UBR] br_10: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [UBR] br_10: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module RetNode2(
  input        clock,
  input        reset,
  output       io_In_enable_ready,
  input        io_In_enable_valid,
  input  [4:0] io_In_enable_bits_taskID,
  input        io_In_enable_bits_control,
  input        io_Out_ready,
  output       io_Out_valid,
  output [4:0] io_Out_bits_enable_taskID,
  output       io_Out_bits_enable_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg  state; // @[RetNode.scala 131:22]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[RetNode.scala 134:31]
  reg [31:0] _RAND_2;
  reg [4:0] output_R_enable_taskID; // @[RetNode.scala 140:25]
  reg [31:0] _RAND_3;
  reg  output_R_enable_control; // @[RetNode.scala 140:25]
  reg [31:0] _RAND_4;
  reg  out_ready_R; // @[RetNode.scala 141:28]
  reg [31:0] _RAND_5;
  reg  out_valid_R; // @[RetNode.scala 142:28]
  reg [31:0] _RAND_6;
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[RetNode.scala 172:23]
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _GEN_8; // @[RetNode.scala 179:28]
  wire  _GEN_9; // @[RetNode.scala 179:28]
  wire  _T_13; // @[RetNode.scala 198:17]
  wire  _T_14; // @[RetNode.scala 198:17]
  wire  _GEN_22; // @[RetNode.scala 198:17]
  wire  _GEN_23; // @[RetNode.scala 198:17]
  wire  _GEN_24; // @[RetNode.scala 198:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_9 = io_In_enable_ready & io_In_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_10 ? 1'h0 : out_valid_R; // @[RetNode.scala 172:23]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _GEN_8 = enable_valid_R | _GEN_5; // @[RetNode.scala 179:28]
  assign _GEN_9 = enable_valid_R | state; // @[RetNode.scala 179:28]
  assign _T_13 = $unsigned(reset); // @[RetNode.scala 198:17]
  assign _T_14 = _T_13 == 1'h0; // @[RetNode.scala 198:17]
  assign io_In_enable_ready = ~ enable_valid_R; // @[RetNode.scala 153:22]
  assign io_Out_valid = out_valid_R; // @[RetNode.scala 170:16]
  assign io_Out_bits_enable_taskID = output_R_enable_taskID; // @[RetNode.scala 169:15]
  assign io_Out_bits_enable_control = output_R_enable_control; // @[RetNode.scala 169:15]
  assign _GEN_22 = _T_11 == 1'h0; // @[RetNode.scala 198:17]
  assign _GEN_23 = _GEN_22 & state; // @[RetNode.scala 198:17]
  assign _GEN_24 = _GEN_23 & out_ready_R; // @[RetNode.scala 198:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  output_R_enable_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  output_R_enable_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_9;
      end else begin
        if (state) begin
          if (out_ready_R) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_9) begin
          enable_valid_R <= io_In_enable_valid;
        end
      end else begin
        if (state) begin
          if (out_ready_R) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_9) begin
              enable_valid_R <= io_In_enable_valid;
            end
          end
        end else begin
          if (_T_9) begin
            enable_valid_R <= io_In_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      output_R_enable_taskID <= 5'h0;
    end else begin
      if (_T_9) begin
        output_R_enable_taskID <= io_In_enable_bits_taskID;
      end
    end
    if (reset) begin
      output_R_enable_control <= 1'h0;
    end else begin
      if (_T_9) begin
        output_R_enable_control <= io_In_enable_bits_control;
      end
    end
    if (reset) begin
      out_ready_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_10) begin
          out_ready_R <= io_Out_ready;
        end
      end else begin
        if (state) begin
          if (out_ready_R) begin
            out_ready_R <= 1'h0;
          end else begin
            if (_T_10) begin
              out_ready_R <= io_Out_ready;
            end
          end
        end else begin
          if (_T_10) begin
            out_ready_R <= io_Out_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        out_valid_R <= _GEN_8;
      end else begin
        if (state) begin
          if (out_ready_R) begin
            out_valid_R <= 1'h0;
          end else begin
            if (_T_10) begin
              out_valid_R <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            out_valid_R <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_24 & _T_14) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [RET] ret_11: Output fired @ %d\n",output_R_enable_taskID,value); // @[RetNode.scala 198:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [31:0] io_Out_2_bits_data,
  input         io_Out_3_ready,
  output        io_Out_3_valid,
  output [31:0] io_Out_3_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_4;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_5;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_6;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_7;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_8;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_9;
  reg  out_valid_R_2; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_10;
  reg  out_valid_R_3; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_11;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_12;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_13;
  reg  fire_R_2; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_14;
  reg  fire_R_3; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_15;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_17; // @[Bitwise.scala 108:18]
  wire  _T_18; // @[Bitwise.scala 108:44]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  _T_22; // @[Decoupled.scala 40:37]
  wire  _GEN_24; // @[PhiNode.scala 258:26]
  wire  _GEN_25; // @[PhiNode.scala 258:26]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _GEN_26; // @[PhiNode.scala 258:26]
  wire  _GEN_27; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  wire  fire_mask_2; // @[PhiNode.scala 265:74]
  wire  fire_mask_3; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_16;
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_29; // @[PhiNode.scala 268:37]
  wire  _T_30; // @[PhiNode.scala 277:27]
  wire  _T_31; // @[PhiNode.scala 283:19]
  wire  _T_32; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_36; // @[PhiNode.scala 283:19]
  wire  _GEN_39; // @[PhiNode.scala 277:46]
  wire  _GEN_40; // @[PhiNode.scala 277:46]
  wire  _GEN_41; // @[PhiNode.scala 277:46]
  wire  _GEN_42; // @[PhiNode.scala 277:46]
  wire  _T_35; // @[Conditional.scala 37:30]
  wire  _T_36; // @[PhiNode.scala 299:31]
  wire  _T_37; // @[PhiNode.scala 299:31]
  wire  _T_38; // @[PhiNode.scala 299:31]
  wire  _T_42; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_80; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_128; // @[Conditional.scala 39:67]
  wire  _GEN_174; // @[PhiNode.scala 283:19]
  wire  _GEN_175; // @[PhiNode.scala 283:19]
  wire  _GEN_177; // @[PhiNode.scala 291:19]
  wire  _GEN_178; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_17 = mask_R[0]; // @[Bitwise.scala 108:18]
  assign _T_18 = mask_R[1]; // @[Bitwise.scala 108:44]
  assign _T_19 = {_T_17,_T_18}; // @[Cat.scala 29:58]
  assign sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  assign _GEN_19 = sel ? in_data_R_1_data : 32'h0; // @[PhiNode.scala 253:20]
  assign _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_20 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = _T_21 | fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign _T_22 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_24 = _T_22 | fire_R_2; // @[PhiNode.scala 258:26]
  assign _GEN_25 = _T_22 ? 1'h0 : out_valid_R_2; // @[PhiNode.scala 258:26]
  assign _T_23 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_26 = _T_23 | fire_R_3; // @[PhiNode.scala 258:26]
  assign _GEN_27 = _T_23 ? 1'h0 : out_valid_R_3; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 265:74]
  assign fire_mask_2 = fire_R_2 | _T_22; // @[PhiNode.scala 265:74]
  assign fire_mask_3 = fire_R_3 | _T_23; // @[PhiNode.scala 265:74]
  assign _T_28 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_29 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_30 = enable_valid_R & _T_29; // @[PhiNode.scala 277:27]
  assign _T_31 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_32 = _T_31 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_36 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_39 = _T_30 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_40 = _T_30 | _GEN_23; // @[PhiNode.scala 277:46]
  assign _GEN_41 = _T_30 | _GEN_25; // @[PhiNode.scala 277:46]
  assign _GEN_42 = _T_30 | _GEN_27; // @[PhiNode.scala 277:46]
  assign _T_35 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_37 = _T_36 & fire_mask_2; // @[PhiNode.scala 299:31]
  assign _T_38 = _T_37 & fire_mask_3; // @[PhiNode.scala 299:31]
  assign _T_42 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_80 = _T_42 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_128 = _T_35 ? _GEN_19 : _GEN_80; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_28 ? _GEN_19 : _GEN_128; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_data = _T_28 ? _GEN_19 : _GEN_128; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_2_valid = out_valid_R_2; // @[PhiNode.scala 254:21]
  assign io_Out_2_bits_data = _T_28 ? _GEN_19 : _GEN_128; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_3_valid = out_valid_R_3; // @[PhiNode.scala 254:21]
  assign io_Out_3_bits_data = _T_28 ? _GEN_19 : _GEN_128; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_174 = _T_28 & _T_30; // @[PhiNode.scala 283:19]
  assign _GEN_175 = _GEN_174 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_177 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_178 = _GEN_174 & _GEN_177; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mask_R = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mask_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fire_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_R_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_R_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  fire_R_3 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  state = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_28) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_28) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_28) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_28) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_28) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_28) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_28) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_28) begin
        out_valid_R_0 <= _GEN_39;
      end else begin
        if (_T_20) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_28) begin
        out_valid_R_1 <= _GEN_40;
      end else begin
        if (_T_21) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_28) begin
        out_valid_R_2 <= _GEN_41;
      end else begin
        if (_T_22) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_28) begin
        out_valid_R_3 <= _GEN_42;
      end else begin
        if (_T_23) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_28) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_28) begin
        fire_R_1 <= _GEN_22;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            fire_R_1 <= 1'h0;
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              fire_R_1 <= 1'h0;
            end else begin
              fire_R_1 <= _GEN_22;
            end
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end
      end
    end
    if (reset) begin
      fire_R_2 <= 1'h0;
    end else begin
      if (_T_28) begin
        fire_R_2 <= _GEN_24;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            fire_R_2 <= 1'h0;
          end else begin
            fire_R_2 <= _GEN_24;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              fire_R_2 <= 1'h0;
            end else begin
              fire_R_2 <= _GEN_24;
            end
          end else begin
            fire_R_2 <= _GEN_24;
          end
        end
      end
    end
    if (reset) begin
      fire_R_3 <= 1'h0;
    end else begin
      if (_T_28) begin
        fire_R_3 <= _GEN_26;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            fire_R_3 <= 1'h0;
          end else begin
            fire_R_3 <= _GEN_26;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              fire_R_3 <= 1'h0;
            end else begin
              fire_R_3 <= _GEN_26;
            end
          end else begin
            fire_R_3 <= _GEN_26;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_28) begin
        if (_T_30) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_32) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [PHI] phi_conv_s1_y_031312: Output fired @ %d, Value: %d\n",_GEN_36,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_178 & _T_32) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [PHI] phi_conv_s1_y_031312: Output flushed @ %d, Value: %d\n",_GEN_36,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_2(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire [18:0] _T_9; // @[Alu.scala 184:47]
  wire [524318:0] _GEN_0; // @[Alu.scala 184:38]
  wire [524318:0] _T_10; // @[Alu.scala 184:38]
  assign _T_9 = io_in2[18:0]; // @[Alu.scala 184:47]
  assign _GEN_0 = {{524287'd0}, io_in1}; // @[Alu.scala 184:38]
  assign _T_10 = _GEN_0 << _T_9; // @[Alu.scala 184:38]
  assign io_out = _T_10[31:0]; // @[Alu.scala 236:10]
endmodule
module ComputeNode_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_2 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul113: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_3(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  assign io_out = io_in1 | io_in2; // @[Alu.scala 236:10]
endmodule
module ComputeNode_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_3 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add214: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul315: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_5(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  assign io_out = io_in1 - io_in2; // @[Alu.scala 236:10]
endmodule
module ComputeNode_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_5 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_sub16: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_6(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h2;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add417: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_7(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul518: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_8(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_5 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_sub619: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_9(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul720: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_10(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h1f;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul821: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UBranchNode_1(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_enable_bits_control,
  input        io_Out_0_ready,
  output       io_Out_0_valid,
  output [4:0] io_Out_0_bits_taskID,
  output       io_Out_0_bits_control
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  state; // @[BranchNode.scala 586:22]
  reg [31:0] _RAND_6;
  wire  _T_11; // @[Conditional.scala 37:30]
  wire  _T_14; // @[HandShaking.scala 652:72]
  wire  _T_15; // @[BranchNode.scala 615:19]
  wire  _T_16; // @[BranchNode.scala 615:19]
  wire  _GEN_6; // @[BranchNode.scala 609:46]
  wire  _GEN_8; // @[BranchNode.scala 609:46]
  wire  _T_22; // @[HandShaking.scala 648:29]
  wire  _GEN_26; // @[BranchNode.scala 615:19]
  wire  _GEN_27; // @[BranchNode.scala 615:19]
  wire  _GEN_29; // @[BranchNode.scala 621:19]
  wire  _GEN_30; // @[BranchNode.scala 621:19]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _T_15 = $unsigned(reset); // @[BranchNode.scala 615:19]
  assign _T_16 = _T_15 == 1'h0; // @[BranchNode.scala 615:19]
  assign _GEN_6 = enable_valid_R | state; // @[BranchNode.scala 609:46]
  assign _GEN_8 = enable_valid_R | out_valid_R_0; // @[BranchNode.scala 609:46]
  assign _T_22 = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = _T_11 ? _GEN_8 : out_valid_R_0; // @[HandShaking.scala 555:21 BranchNode.scala 612:32]
  assign io_Out_0_bits_taskID = enable_R_taskID; // @[BranchNode.scala 605:25]
  assign io_Out_0_bits_control = enable_R_control; // @[BranchNode.scala 605:25]
  assign _GEN_26 = _T_11 & enable_valid_R; // @[BranchNode.scala 615:19]
  assign _GEN_27 = _GEN_26 & enable_R_control; // @[BranchNode.scala 615:19]
  assign _GEN_29 = enable_R_control == 1'h0; // @[BranchNode.scala 621:19]
  assign _GEN_30 = _GEN_26 & _GEN_29; // @[BranchNode.scala 621:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_6) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_6) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_11) begin
        if (enable_valid_R) begin
          out_valid_R_0 <= _T_14;
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_11) begin
        state <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_27 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [UBR] br_22: Output fired [T] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 615:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_30 & _T_16) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [UBR] br_22: Output fired [F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 621:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_11(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_inc12023: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UALU_12(
  input  [31:0] io_in1,
  input  [31:0] io_in2,
  output [31:0] io_out
);
  wire  _T_21; // @[Alu.scala 190:38]
  assign _T_21 = io_in1 == io_in2; // @[Alu.scala 190:38]
  assign io_out = {{31'd0}, _T_21}; // @[Alu.scala 236:10]
endmodule
module ComputeNode_12(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_12 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h1f;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] icmp_exitcond31424: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_8;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_9;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_10;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_12;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_13;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_14;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CBR] br_25: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CBR] br_25: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module PhiFastNode_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input         io_enable_bits_control,
  output        io_InData_0_ready,
  input         io_InData_0_valid,
  input  [4:0]  io_InData_0_bits_taskID,
  output        io_InData_1_ready,
  input         io_InData_1_valid,
  input  [4:0]  io_InData_1_bits_taskID,
  input  [31:0] io_InData_1_bits_data,
  output        io_Mask_ready,
  input         io_Mask_valid,
  input  [1:0]  io_Mask_bits,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [31:0] io_Out_2_bits_data,
  input         io_Out_3_ready,
  output        io_Out_3_valid,
  output [31:0] io_Out_3_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] in_data_R_1_data; // @[PhiNode.scala 197:26]
  reg [31:0] _RAND_1;
  reg  in_data_valid_R_0; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_2;
  reg  in_data_valid_R_1; // @[PhiNode.scala 198:32]
  reg [31:0] _RAND_3;
  reg  enable_R_control; // @[PhiNode.scala 201:25]
  reg [31:0] _RAND_4;
  reg  enable_valid_R; // @[PhiNode.scala 202:31]
  reg [31:0] _RAND_5;
  reg [1:0] mask_R; // @[PhiNode.scala 205:23]
  reg [31:0] _RAND_6;
  reg  mask_valid_R; // @[PhiNode.scala 206:29]
  reg [31:0] _RAND_7;
  reg  out_valid_R_0; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_8;
  reg  out_valid_R_1; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_9;
  reg  out_valid_R_2; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_10;
  reg  out_valid_R_3; // @[PhiNode.scala 209:49]
  reg [31:0] _RAND_11;
  reg  fire_R_0; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_12;
  reg  fire_R_1; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_13;
  reg  fire_R_2; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_14;
  reg  fire_R_3; // @[PhiNode.scala 211:44]
  reg [31:0] _RAND_15;
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_2; // @[PhiNode.scala 215:24]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_5; // @[PhiNode.scala 222:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[PhiNode.scala 230:29]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[PhiNode.scala 230:29]
  wire  _T_17; // @[Bitwise.scala 108:18]
  wire  _T_18; // @[Bitwise.scala 108:44]
  wire [1:0] _T_19; // @[Cat.scala 29:58]
  wire  sel; // @[CircuitMath.scala 30:8]
  wire [31:0] _GEN_19; // @[PhiNode.scala 253:20]
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_20; // @[PhiNode.scala 258:26]
  wire  _GEN_21; // @[PhiNode.scala 258:26]
  wire  _T_21; // @[Decoupled.scala 40:37]
  wire  _GEN_22; // @[PhiNode.scala 258:26]
  wire  _GEN_23; // @[PhiNode.scala 258:26]
  wire  _T_22; // @[Decoupled.scala 40:37]
  wire  _GEN_24; // @[PhiNode.scala 258:26]
  wire  _GEN_25; // @[PhiNode.scala 258:26]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _GEN_26; // @[PhiNode.scala 258:26]
  wire  _GEN_27; // @[PhiNode.scala 258:26]
  wire  fire_mask_0; // @[PhiNode.scala 265:74]
  wire  fire_mask_1; // @[PhiNode.scala 265:74]
  wire  fire_mask_2; // @[PhiNode.scala 265:74]
  wire  fire_mask_3; // @[PhiNode.scala 265:74]
  reg [1:0] state; // @[PhiNode.scala 273:22]
  reg [31:0] _RAND_16;
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_29; // @[PhiNode.scala 268:37]
  wire  _T_30; // @[PhiNode.scala 277:27]
  wire  _T_31; // @[PhiNode.scala 283:19]
  wire  _T_32; // @[PhiNode.scala 283:19]
  wire [4:0] _GEN_36; // @[PhiNode.scala 283:19]
  wire  _GEN_39; // @[PhiNode.scala 277:46]
  wire  _GEN_40; // @[PhiNode.scala 277:46]
  wire  _GEN_41; // @[PhiNode.scala 277:46]
  wire  _GEN_42; // @[PhiNode.scala 277:46]
  wire  _T_35; // @[Conditional.scala 37:30]
  wire  _T_36; // @[PhiNode.scala 299:31]
  wire  _T_37; // @[PhiNode.scala 299:31]
  wire  _T_38; // @[PhiNode.scala 299:31]
  wire  _T_42; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_80; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_128; // @[Conditional.scala 39:67]
  wire  _GEN_174; // @[PhiNode.scala 283:19]
  wire  _GEN_175; // @[PhiNode.scala 283:19]
  wire  _GEN_177; // @[PhiNode.scala 291:19]
  wire  _GEN_178; // @[PhiNode.scala 291:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_10 = io_Mask_ready & io_Mask_valid; // @[Decoupled.scala 40:37]
  assign _GEN_2 = _T_10 | mask_valid_R; // @[PhiNode.scala 215:24]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_5 = _T_12 | enable_valid_R; // @[PhiNode.scala 222:26]
  assign _T_14 = io_InData_0_ready & io_InData_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | in_data_valid_R_0; // @[PhiNode.scala 230:29]
  assign _T_16 = io_InData_1_ready & io_InData_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_16 | in_data_valid_R_1; // @[PhiNode.scala 230:29]
  assign _T_17 = mask_R[0]; // @[Bitwise.scala 108:18]
  assign _T_18 = mask_R[1]; // @[Bitwise.scala 108:44]
  assign _T_19 = {_T_17,_T_18}; // @[Cat.scala 29:58]
  assign sel = _T_19[1]; // @[CircuitMath.scala 30:8]
  assign _GEN_19 = sel ? in_data_R_1_data : 32'h0; // @[PhiNode.scala 253:20]
  assign _T_20 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_20 = _T_20 | fire_R_0; // @[PhiNode.scala 258:26]
  assign _GEN_21 = _T_20 ? 1'h0 : out_valid_R_0; // @[PhiNode.scala 258:26]
  assign _T_21 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _GEN_22 = _T_21 | fire_R_1; // @[PhiNode.scala 258:26]
  assign _GEN_23 = _T_21 ? 1'h0 : out_valid_R_1; // @[PhiNode.scala 258:26]
  assign _T_22 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _GEN_24 = _T_22 | fire_R_2; // @[PhiNode.scala 258:26]
  assign _GEN_25 = _T_22 ? 1'h0 : out_valid_R_2; // @[PhiNode.scala 258:26]
  assign _T_23 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _GEN_26 = _T_23 | fire_R_3; // @[PhiNode.scala 258:26]
  assign _GEN_27 = _T_23 ? 1'h0 : out_valid_R_3; // @[PhiNode.scala 258:26]
  assign fire_mask_0 = fire_R_0 | _T_20; // @[PhiNode.scala 265:74]
  assign fire_mask_1 = fire_R_1 | _T_21; // @[PhiNode.scala 265:74]
  assign fire_mask_2 = fire_R_2 | _T_22; // @[PhiNode.scala 265:74]
  assign fire_mask_3 = fire_R_3 | _T_23; // @[PhiNode.scala 265:74]
  assign _T_28 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_29 = in_data_valid_R_0 & in_data_valid_R_1; // @[PhiNode.scala 268:37]
  assign _T_30 = enable_valid_R & _T_29; // @[PhiNode.scala 277:27]
  assign _T_31 = $unsigned(reset); // @[PhiNode.scala 283:19]
  assign _T_32 = _T_31 == 1'h0; // @[PhiNode.scala 283:19]
  assign _GEN_36 = sel ? io_InData_1_bits_taskID : io_InData_0_bits_taskID; // @[PhiNode.scala 283:19]
  assign _GEN_39 = _T_30 | _GEN_21; // @[PhiNode.scala 277:46]
  assign _GEN_40 = _T_30 | _GEN_23; // @[PhiNode.scala 277:46]
  assign _GEN_41 = _T_30 | _GEN_25; // @[PhiNode.scala 277:46]
  assign _GEN_42 = _T_30 | _GEN_27; // @[PhiNode.scala 277:46]
  assign _T_35 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = fire_mask_0 & fire_mask_1; // @[PhiNode.scala 299:31]
  assign _T_37 = _T_36 & fire_mask_2; // @[PhiNode.scala 299:31]
  assign _T_38 = _T_37 & fire_mask_3; // @[PhiNode.scala 299:31]
  assign _T_42 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _GEN_80 = _T_42 ? 32'h0 : _GEN_19; // @[Conditional.scala 39:67]
  assign _GEN_128 = _T_35 ? _GEN_19 : _GEN_80; // @[Conditional.scala 39:67]
  assign io_enable_ready = ~ enable_valid_R; // @[PhiNode.scala 221:19]
  assign io_InData_0_ready = ~ in_data_valid_R_0; // @[PhiNode.scala 229:24]
  assign io_InData_1_ready = ~ in_data_valid_R_1; // @[PhiNode.scala 229:24]
  assign io_Mask_ready = ~ mask_valid_R; // @[PhiNode.scala 214:17]
  assign io_Out_0_valid = out_valid_R_0; // @[PhiNode.scala 254:21]
  assign io_Out_0_bits_data = _T_28 ? _GEN_19 : _GEN_128; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_1_valid = out_valid_R_1; // @[PhiNode.scala 254:21]
  assign io_Out_1_bits_data = _T_28 ? _GEN_19 : _GEN_128; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_2_valid = out_valid_R_2; // @[PhiNode.scala 254:21]
  assign io_Out_2_bits_data = _T_28 ? _GEN_19 : _GEN_128; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign io_Out_3_valid = out_valid_R_3; // @[PhiNode.scala 254:21]
  assign io_Out_3_bits_data = _T_28 ? _GEN_19 : _GEN_128; // @[PhiNode.scala 253:20 PhiNode.scala 325:42]
  assign _GEN_174 = _T_28 & _T_30; // @[PhiNode.scala 283:19]
  assign _GEN_175 = _GEN_174 & enable_R_control; // @[PhiNode.scala 283:19]
  assign _GEN_177 = enable_R_control == 1'h0; // @[PhiNode.scala 291:19]
  assign _GEN_178 = _GEN_174 & _GEN_177; // @[PhiNode.scala 291:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  in_data_R_1_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  in_data_valid_R_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  in_data_valid_R_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_control = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_valid_R = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mask_R = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mask_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  fire_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_R_1 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  fire_R_2 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  fire_R_3 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  state = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      in_data_R_1_data <= 32'h0;
    end else begin
      if (_T_28) begin
        if (_T_16) begin
          in_data_R_1_data <= io_InData_1_bits_data;
        end
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            in_data_R_1_data <= 32'h0;
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              in_data_R_1_data <= 32'h0;
            end else begin
              if (_T_16) begin
                in_data_R_1_data <= io_InData_1_bits_data;
              end
            end
          end else begin
            if (_T_16) begin
              in_data_R_1_data <= io_InData_1_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_0 <= 1'h0;
    end else begin
      if (_T_28) begin
        in_data_valid_R_0 <= _GEN_9;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            in_data_valid_R_0 <= 1'h0;
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              in_data_valid_R_0 <= 1'h0;
            end else begin
              in_data_valid_R_0 <= _GEN_9;
            end
          end else begin
            in_data_valid_R_0 <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      in_data_valid_R_1 <= 1'h0;
    end else begin
      if (_T_28) begin
        in_data_valid_R_1 <= _GEN_13;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            in_data_valid_R_1 <= 1'h0;
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              in_data_valid_R_1 <= 1'h0;
            end else begin
              in_data_valid_R_1 <= _GEN_13;
            end
          end else begin
            in_data_valid_R_1 <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_28) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              enable_R_control <= 1'h0;
            end else begin
              if (_T_12) begin
                enable_R_control <= io_enable_bits_control;
              end
            end
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_28) begin
        enable_valid_R <= _GEN_5;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              enable_valid_R <= 1'h0;
            end else begin
              enable_valid_R <= _GEN_5;
            end
          end else begin
            enable_valid_R <= _GEN_5;
          end
        end
      end
    end
    if (reset) begin
      mask_R <= 2'h0;
    end else begin
      if (_T_28) begin
        if (_T_10) begin
          mask_R <= io_Mask_bits;
        end
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            mask_R <= 2'h0;
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              mask_R <= 2'h0;
            end else begin
              if (_T_10) begin
                mask_R <= io_Mask_bits;
              end
            end
          end else begin
            if (_T_10) begin
              mask_R <= io_Mask_bits;
            end
          end
        end
      end
    end
    if (reset) begin
      mask_valid_R <= 1'h0;
    end else begin
      if (_T_28) begin
        mask_valid_R <= _GEN_2;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            mask_valid_R <= 1'h0;
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              mask_valid_R <= 1'h0;
            end else begin
              mask_valid_R <= _GEN_2;
            end
          end else begin
            mask_valid_R <= _GEN_2;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_28) begin
        out_valid_R_0 <= _GEN_39;
      end else begin
        if (_T_20) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_28) begin
        out_valid_R_1 <= _GEN_40;
      end else begin
        if (_T_21) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_28) begin
        out_valid_R_2 <= _GEN_41;
      end else begin
        if (_T_22) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_28) begin
        out_valid_R_3 <= _GEN_42;
      end else begin
        if (_T_23) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_28) begin
        fire_R_0 <= _GEN_20;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              fire_R_0 <= 1'h0;
            end else begin
              fire_R_0 <= _GEN_20;
            end
          end else begin
            fire_R_0 <= _GEN_20;
          end
        end
      end
    end
    if (reset) begin
      fire_R_1 <= 1'h0;
    end else begin
      if (_T_28) begin
        fire_R_1 <= _GEN_22;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            fire_R_1 <= 1'h0;
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              fire_R_1 <= 1'h0;
            end else begin
              fire_R_1 <= _GEN_22;
            end
          end else begin
            fire_R_1 <= _GEN_22;
          end
        end
      end
    end
    if (reset) begin
      fire_R_2 <= 1'h0;
    end else begin
      if (_T_28) begin
        fire_R_2 <= _GEN_24;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            fire_R_2 <= 1'h0;
          end else begin
            fire_R_2 <= _GEN_24;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              fire_R_2 <= 1'h0;
            end else begin
              fire_R_2 <= _GEN_24;
            end
          end else begin
            fire_R_2 <= _GEN_24;
          end
        end
      end
    end
    if (reset) begin
      fire_R_3 <= 1'h0;
    end else begin
      if (_T_28) begin
        fire_R_3 <= _GEN_26;
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            fire_R_3 <= 1'h0;
          end else begin
            fire_R_3 <= _GEN_26;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              fire_R_3 <= 1'h0;
            end else begin
              fire_R_3 <= _GEN_26;
            end
          end else begin
            fire_R_3 <= _GEN_26;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_28) begin
        if (_T_30) begin
          if (enable_R_control) begin
            state <= 2'h1;
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_35) begin
          if (_T_38) begin
            state <= 2'h0;
          end
        end else begin
          if (_T_42) begin
            if (_T_38) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_175 & _T_32) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [PHI] phi_conv_s1_x_031226: Output fired @ %d, Value: %d\n",_GEN_36,value,_GEN_19); // @[PhiNode.scala 283:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_178 & _T_32) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [PHI] phi_conv_s1_x_031226: Output flushed @ %d, Value: %d\n",_GEN_36,value,_GEN_19); // @[PhiNode.scala 291:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_13(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add1327: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_8(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [4:0]  io_Out_1_bits_taskID,
  output [31:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [4:0]  io_Out_2_bits_taskID,
  output [31:0] io_Out_2_bits_data,
  input         io_Out_3_ready,
  output        io_Out_3_valid,
  output [4:0]  io_Out_3_bits_taskID,
  output [31:0] io_Out_3_bits_data,
  input         io_Out_4_ready,
  output        io_Out_4_valid,
  output [4:0]  io_Out_4_bits_taskID,
  output [31:0] io_Out_4_bits_data,
  input         io_Out_5_ready,
  output        io_Out_5_valid,
  output [4:0]  io_Out_5_bits_taskID,
  output [31:0] io_Out_5_bits_data,
  input         io_Out_6_ready,
  output        io_Out_6_valid,
  output [4:0]  io_Out_6_bits_taskID,
  output [31:0] io_Out_6_bits_data,
  input         io_Out_7_ready,
  output        io_Out_7_valid,
  output [4:0]  io_Out_7_bits_taskID,
  output [31:0] io_Out_7_bits_data,
  input         io_Out_8_ready,
  output        io_Out_8_valid,
  output [4:0]  io_Out_8_bits_taskID,
  output [31:0] io_Out_8_bits_data,
  input         io_Out_9_ready,
  output        io_Out_9_valid,
  output [4:0]  io_Out_9_bits_taskID,
  output [31:0] io_Out_9_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_ready_R_2; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_5;
  reg  out_ready_R_3; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_6;
  reg  out_ready_R_4; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_7;
  reg  out_ready_R_5; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_8;
  reg  out_ready_R_6; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_9;
  reg  out_ready_R_7; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_10;
  reg  out_ready_R_8; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_11;
  reg  out_ready_R_9; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_12;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_13;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_14;
  reg  out_valid_R_2; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_15;
  reg  out_valid_R_3; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_16;
  reg  out_valid_R_4; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_17;
  reg  out_valid_R_5; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_18;
  reg  out_valid_R_6; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_19;
  reg  out_valid_R_7; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_20;
  reg  out_valid_R_8; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_21;
  reg  out_valid_R_9; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_22;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_5; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _T_12; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_23;
  wire [14:0] _T_15; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_24;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_25;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_26;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_27;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_28;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_29;
  wire  _T_20; // @[Decoupled.scala 40:37]
  wire  _GEN_27; // @[GepNode.scala 905:31]
  wire  _T_22; // @[Decoupled.scala 40:37]
  wire  _GEN_31; // @[GepNode.scala 912:28]
  wire [34:0] seek_value; // @[GepNode.scala 920:21]
  wire [34:0] _GEN_113; // @[GepNode.scala 928:35]
  wire [34:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_24; // @[Conditional.scala 37:30]
  wire  _T_25; // @[GepNode.scala 944:27]
  wire  _T_26; // @[GepNode.scala 944:48]
  wire  _T_37; // @[HandShaking.scala 232:72]
  wire  _T_38; // @[HandShaking.scala 232:72]
  wire  _T_39; // @[HandShaking.scala 232:72]
  wire  _T_40; // @[HandShaking.scala 232:72]
  wire  _T_41; // @[HandShaking.scala 232:72]
  wire  _T_42; // @[HandShaking.scala 232:72]
  wire  _T_43; // @[HandShaking.scala 232:72]
  wire  _T_44; // @[HandShaking.scala 232:72]
  wire  _T_45; // @[HandShaking.scala 232:72]
  wire  _T_46; // @[HandShaking.scala 232:72]
  wire  _GEN_42; // @[GepNode.scala 944:78]
  wire  _T_58; // @[HandShaking.scala 217:83]
  wire  _T_59; // @[HandShaking.scala 217:83]
  wire  _T_60; // @[HandShaking.scala 217:83]
  wire  _T_61; // @[HandShaking.scala 217:83]
  wire  _T_62; // @[HandShaking.scala 217:83]
  wire  _T_63; // @[HandShaking.scala 217:83]
  wire  _T_64; // @[HandShaking.scala 217:83]
  wire  _T_65; // @[HandShaking.scala 217:83]
  wire  _T_66; // @[HandShaking.scala 217:83]
  wire  _T_67; // @[HandShaking.scala 217:83]
  wire  _T_68; // @[HandShaking.scala 218:27]
  wire  _T_69; // @[HandShaking.scala 218:27]
  wire  _T_70; // @[HandShaking.scala 218:27]
  wire  _T_71; // @[HandShaking.scala 218:27]
  wire  _T_72; // @[HandShaking.scala 218:27]
  wire  _T_73; // @[HandShaking.scala 218:27]
  wire  _T_74; // @[HandShaking.scala 218:27]
  wire  _T_75; // @[HandShaking.scala 218:27]
  wire  _T_76; // @[HandShaking.scala 218:27]
  wire  _T_79; // @[GepNode.scala 964:17]
  wire  _T_80; // @[GepNode.scala 964:17]
  wire  _GEN_114; // @[GepNode.scala 964:17]
  wire  _GEN_115; // @[GepNode.scala 964:17]
  wire  _GEN_116; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_Out_3_ready & io_Out_3_valid; // @[Decoupled.scala 40:37]
  assign _T_5 = io_Out_4_ready & io_Out_4_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_Out_5_ready & io_Out_5_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = io_Out_6_ready & io_Out_6_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = io_Out_7_ready & io_Out_7_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_8_ready & io_Out_8_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_Out_9_ready & io_Out_9_valid; // @[Decoupled.scala 40:37]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_15 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_20 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_27 = _T_20 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_22 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_31 = _T_22 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h4; // @[GepNode.scala 920:21]
  assign _GEN_113 = {{3'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_113 + seek_value; // @[GepNode.scala 928:35]
  assign _T_24 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_25 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_26 = _T_25 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_37 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_38 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_39 = _T_3 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_40 = _T_4 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_41 = _T_5 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_42 = _T_6 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_43 = _T_7 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_44 = _T_8 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_45 = _T_9 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_46 = _T_10 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_42 = _T_26 | state; // @[GepNode.scala 944:78]
  assign _T_58 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_59 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_60 = out_ready_R_2 | _T_3; // @[HandShaking.scala 217:83]
  assign _T_61 = out_ready_R_3 | _T_4; // @[HandShaking.scala 217:83]
  assign _T_62 = out_ready_R_4 | _T_5; // @[HandShaking.scala 217:83]
  assign _T_63 = out_ready_R_5 | _T_6; // @[HandShaking.scala 217:83]
  assign _T_64 = out_ready_R_6 | _T_7; // @[HandShaking.scala 217:83]
  assign _T_65 = out_ready_R_7 | _T_8; // @[HandShaking.scala 217:83]
  assign _T_66 = out_ready_R_8 | _T_9; // @[HandShaking.scala 217:83]
  assign _T_67 = out_ready_R_9 | _T_10; // @[HandShaking.scala 217:83]
  assign _T_68 = _T_58 & _T_59; // @[HandShaking.scala 218:27]
  assign _T_69 = _T_68 & _T_60; // @[HandShaking.scala 218:27]
  assign _T_70 = _T_69 & _T_61; // @[HandShaking.scala 218:27]
  assign _T_71 = _T_70 & _T_62; // @[HandShaking.scala 218:27]
  assign _T_72 = _T_71 & _T_63; // @[HandShaking.scala 218:27]
  assign _T_73 = _T_72 & _T_64; // @[HandShaking.scala 218:27]
  assign _T_74 = _T_73 & _T_65; // @[HandShaking.scala 218:27]
  assign _T_75 = _T_74 & _T_66; // @[HandShaking.scala 218:27]
  assign _T_76 = _T_75 & _T_67; // @[HandShaking.scala 218:27]
  assign _T_79 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_80 = _T_79 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_Out_1_valid = out_valid_R_1; // @[HandShaking.scala 180:21]
  assign io_Out_1_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_1_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_Out_2_valid = out_valid_R_2; // @[HandShaking.scala 180:21]
  assign io_Out_2_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_2_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_Out_3_valid = out_valid_R_3; // @[HandShaking.scala 180:21]
  assign io_Out_3_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_3_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_Out_4_valid = out_valid_R_4; // @[HandShaking.scala 180:21]
  assign io_Out_4_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_4_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_Out_5_valid = out_valid_R_5; // @[HandShaking.scala 180:21]
  assign io_Out_5_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_5_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_Out_6_valid = out_valid_R_6; // @[HandShaking.scala 180:21]
  assign io_Out_6_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_6_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_Out_7_valid = out_valid_R_7; // @[HandShaking.scala 180:21]
  assign io_Out_7_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_7_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_Out_8_valid = out_valid_R_8; // @[HandShaking.scala 180:21]
  assign io_Out_8_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_8_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_Out_9_valid = out_valid_R_9; // @[HandShaking.scala 180:21]
  assign io_Out_9_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_9_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_114 = _T_24 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_115 = _GEN_114 & state; // @[GepNode.scala 964:17]
  assign _GEN_116 = _GEN_115 & _T_76; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_ready_R_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_ready_R_4 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_ready_R_5 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  out_ready_R_6 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  out_ready_R_7 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_ready_R_8 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  out_ready_R_9 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  out_valid_R_3 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  out_valid_R_4 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  out_valid_R_5 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  out_valid_R_6 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  out_valid_R_7 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  out_valid_R_8 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  out_valid_R_9 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  value = _RAND_23[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_24[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  base_addr_R_data = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  idx_R_0_data = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  state = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_12) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_12) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_3) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_4) begin
          out_ready_R_3 <= io_Out_3_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_3 <= 1'h0;
          end else begin
            if (_T_4) begin
              out_ready_R_3 <= io_Out_3_ready;
            end
          end
        end else begin
          if (_T_4) begin
            out_ready_R_3 <= io_Out_3_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_4 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_5) begin
          out_ready_R_4 <= io_Out_4_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_4 <= 1'h0;
          end else begin
            if (_T_5) begin
              out_ready_R_4 <= io_Out_4_ready;
            end
          end
        end else begin
          if (_T_5) begin
            out_ready_R_4 <= io_Out_4_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_5 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_6) begin
          out_ready_R_5 <= io_Out_5_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_5 <= 1'h0;
          end else begin
            if (_T_6) begin
              out_ready_R_5 <= io_Out_5_ready;
            end
          end
        end else begin
          if (_T_6) begin
            out_ready_R_5 <= io_Out_5_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_6 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_7) begin
          out_ready_R_6 <= io_Out_6_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_6 <= 1'h0;
          end else begin
            if (_T_7) begin
              out_ready_R_6 <= io_Out_6_ready;
            end
          end
        end else begin
          if (_T_7) begin
            out_ready_R_6 <= io_Out_6_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_7 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_8) begin
          out_ready_R_7 <= io_Out_7_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_7 <= 1'h0;
          end else begin
            if (_T_8) begin
              out_ready_R_7 <= io_Out_7_ready;
            end
          end
        end else begin
          if (_T_8) begin
            out_ready_R_7 <= io_Out_7_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_8 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_9) begin
          out_ready_R_8 <= io_Out_8_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_8 <= 1'h0;
          end else begin
            if (_T_9) begin
              out_ready_R_8 <= io_Out_8_ready;
            end
          end
        end else begin
          if (_T_9) begin
            out_ready_R_8 <= io_Out_8_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_9 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_10) begin
          out_ready_R_9 <= io_Out_9_ready;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            out_ready_R_9 <= 1'h0;
          end else begin
            if (_T_10) begin
              out_ready_R_9 <= io_Out_9_ready;
            end
          end
        end else begin
          if (_T_10) begin
            out_ready_R_9 <= io_Out_9_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_0 <= _T_37;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_1 <= _T_38;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_2 <= _T_39;
        end else begin
          if (_T_3) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_3) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_3 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_3 <= _T_40;
        end else begin
          if (_T_4) begin
            out_valid_R_3 <= 1'h0;
          end
        end
      end else begin
        if (_T_4) begin
          out_valid_R_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_4 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_4 <= _T_41;
        end else begin
          if (_T_5) begin
            out_valid_R_4 <= 1'h0;
          end
        end
      end else begin
        if (_T_5) begin
          out_valid_R_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_5 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_5 <= _T_42;
        end else begin
          if (_T_6) begin
            out_valid_R_5 <= 1'h0;
          end
        end
      end else begin
        if (_T_6) begin
          out_valid_R_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_6 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_6 <= _T_43;
        end else begin
          if (_T_7) begin
            out_valid_R_6 <= 1'h0;
          end
        end
      end else begin
        if (_T_7) begin
          out_valid_R_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_7 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_7 <= _T_44;
        end else begin
          if (_T_8) begin
            out_valid_R_7 <= 1'h0;
          end
        end
      end else begin
        if (_T_8) begin
          out_valid_R_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_8 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_8 <= _T_45;
        end else begin
          if (_T_9) begin
            out_valid_R_8 <= 1'h0;
          end
        end
      end else begin
        if (_T_9) begin
          out_valid_R_8 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_9 <= 1'h0;
    end else begin
      if (_T_24) begin
        if (_T_26) begin
          out_valid_R_9 <= _T_46;
        end else begin
          if (_T_10) begin
            out_valid_R_9 <= 1'h0;
          end
        end
      end else begin
        if (_T_10) begin
          out_valid_R_9 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_15;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_24) begin
        if (_T_20) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_20) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_20) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_24) begin
        if (_T_20) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_20) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_20) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_24) begin
        base_addr_valid_R <= _GEN_27;
      end else begin
        if (state) begin
          if (_T_76) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_27;
          end
        end else begin
          base_addr_valid_R <= _GEN_27;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_24) begin
        if (_T_22) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_76) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_22) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_22) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_24) begin
        idx_valid_R_0 <= _GEN_31;
      end else begin
        if (state) begin
          if (_T_76) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_31;
          end
        end else begin
          idx_valid_R_0 <= _GEN_31;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_24) begin
        state <= _GEN_42;
      end else begin
        if (state) begin
          if (_T_76) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_116 & _T_80) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx28: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_29: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_29: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_29: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_30: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_30: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_30: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_14(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add1531: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_15(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_2 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul1632: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_16(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [31:0] io_Out_2_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_ready_R_2; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_7;
  reg  out_valid_R_2; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _T_5; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_9;
  wire [14:0] _T_8; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_10;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_11;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_12;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_13;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_14;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_15;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 74:26]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[ComputeNode.scala 80:27]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[ComputeNode.scala 99:27]
  wire  _T_22; // @[ComputeNode.scala 99:43]
  wire  _T_29; // @[HandShaking.scala 232:72]
  wire  _T_30; // @[HandShaking.scala 232:72]
  wire  _T_31; // @[HandShaking.scala 232:72]
  wire  _T_32; // @[ComputeNode.scala 107:17]
  wire  _T_33; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_23_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_18; // @[ComputeNode.scala 99:61]
  wire  _GEN_27; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _GEN_29; // @[ComputeNode.scala 99:61]
  wire  _GEN_35; // @[ComputeNode.scala 99:61]
  wire  _T_38; // @[HandShaking.scala 217:83]
  wire  _T_39; // @[HandShaking.scala 217:83]
  wire  _T_40; // @[HandShaking.scala 217:83]
  wire  _T_41; // @[HandShaking.scala 218:27]
  wire  _T_42; // @[HandShaking.scala 218:27]
  wire  _GEN_71; // @[ComputeNode.scala 107:17]
  UALU_5 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _T_5 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_14 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_16 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_16 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_20 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_22 = _T_21 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_29 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_30 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_31 = _T_3 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_32 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_33 = _T_32 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_23_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_18 = _T_22 ? _T_23_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_27 = _T_22 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_22 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_29 = _T_22 | out_valid_R_2; // @[ComputeNode.scala 99:61]
  assign _GEN_35 = _T_22 | state; // @[ComputeNode.scala 99:61]
  assign _T_38 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_39 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_40 = out_ready_R_2 | _T_3; // @[HandShaking.scala 217:83]
  assign _T_41 = _T_38 & _T_39; // @[HandShaking.scala 218:27]
  assign _T_42 = _T_41 & _T_40; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_20 ? _GEN_27 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_20 ? _GEN_18 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_20 ? _GEN_28 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_20 ? _GEN_18 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_2_valid = _T_20 ? _GEN_29 : out_valid_R_2; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_2_bits_data = _T_20 ? _GEN_18 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_71 = _T_20 & _T_22; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value = _RAND_9[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  left_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  left_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  right_R_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  right_valid_R = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_data_R = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_5) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_5) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_5) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_5) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_5) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_3) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          out_valid_R_0 <= _T_29;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          out_valid_R_1 <= _T_30;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          out_valid_R_2 <= _T_31;
        end else begin
          if (_T_3) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_3) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_8;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_13;
        end
      end else begin
        left_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_16) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_17;
        end
      end else begin
        right_valid_R <= _GEN_17;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_20) begin
        state <= _GEN_35;
      end else begin
        if (state) begin
          if (_T_42) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_20) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & _T_33) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_sub1733: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_9(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx1834: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_35: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_35: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_35: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ZextNode(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[ZextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[ZextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[ZextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[ZextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[ZextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[ZextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[ZextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[ZextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[ZextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[ZextNode.scala 84:26]
  wire  _GEN_9; // @[ZextNode.scala 84:26]
  wire  fire_mask_0; // @[ZextNode.scala 90:74]
  reg  state; // @[ZextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[ZextNode.scala 93:27]
  wire  _T_16; // @[ZextNode.scala 97:26]
  wire  _T_17; // @[ZextNode.scala 110:28]
  wire  _T_18; // @[ZextNode.scala 117:17]
  wire  _T_19; // @[ZextNode.scala 117:17]
  wire  _GEN_10; // @[ZextNode.scala 110:47]
  wire  _GEN_11; // @[ZextNode.scala 110:47]
  wire  _GEN_42; // @[ZextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ZextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[ZextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[ZextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[ZextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[ZextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[ZextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[ZextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[ZextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[ZextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[ZextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[ZextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[ZextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[ZextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[ZextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[ZextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[ZextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[ZextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[ZextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] sextconv1936: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[ZextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_17(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul2037: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_18(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add2138: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [STORE]st_39: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_40: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_40: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_40: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_19(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add2941: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_10(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx3042: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_43: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_43: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_43: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ZextNode_1(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[ZextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[ZextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[ZextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[ZextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[ZextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[ZextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[ZextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[ZextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[ZextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[ZextNode.scala 84:26]
  wire  _GEN_9; // @[ZextNode.scala 84:26]
  wire  fire_mask_0; // @[ZextNode.scala 90:74]
  reg  state; // @[ZextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[ZextNode.scala 93:27]
  wire  _T_16; // @[ZextNode.scala 97:26]
  wire  _T_17; // @[ZextNode.scala 110:28]
  wire  _T_18; // @[ZextNode.scala 117:17]
  wire  _T_19; // @[ZextNode.scala 117:17]
  wire  _GEN_10; // @[ZextNode.scala 110:47]
  wire  _GEN_11; // @[ZextNode.scala 110:47]
  wire  _GEN_42; // @[ZextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ZextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[ZextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[ZextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[ZextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[ZextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[ZextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[ZextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[ZextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[ZextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[ZextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[ZextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[ZextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[ZextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[ZextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[ZextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[ZextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[ZextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[ZextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] sextconv3244: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[ZextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_20(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul3345: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_21(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add3446: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [STORE]st_47: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_48: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_48: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_48: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_22(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h2;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add4249: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_11(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx4350: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_6(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_51: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_51: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_51: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ZextNode_2(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[ZextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[ZextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[ZextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[ZextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[ZextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[ZextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[ZextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[ZextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[ZextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[ZextNode.scala 84:26]
  wire  _GEN_9; // @[ZextNode.scala 84:26]
  wire  fire_mask_0; // @[ZextNode.scala 90:74]
  reg  state; // @[ZextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[ZextNode.scala 93:27]
  wire  _T_16; // @[ZextNode.scala 97:26]
  wire  _T_17; // @[ZextNode.scala 110:28]
  wire  _T_18; // @[ZextNode.scala 117:17]
  wire  _T_19; // @[ZextNode.scala 117:17]
  wire  _GEN_10; // @[ZextNode.scala 110:47]
  wire  _GEN_11; // @[ZextNode.scala 110:47]
  wire  _GEN_42; // @[ZextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ZextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[ZextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[ZextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[ZextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[ZextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[ZextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[ZextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[ZextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[ZextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[ZextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[ZextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[ZextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[ZextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[ZextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[ZextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[ZextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[ZextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[ZextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] sextconv4552: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[ZextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_23(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul4653: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_24(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add4754: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore_2(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [STORE]st_55: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_7(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_56: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_56: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_56: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_25(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_2 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul5257: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_26(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [31:0] io_Out_2_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_ready_R_2; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_7;
  reg  out_valid_R_2; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _T_5; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_9;
  wire [14:0] _T_8; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_10;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_11;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_12;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_13;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_14;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_15;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 74:26]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[ComputeNode.scala 80:27]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[ComputeNode.scala 99:27]
  wire  _T_22; // @[ComputeNode.scala 99:43]
  wire  _T_29; // @[HandShaking.scala 232:72]
  wire  _T_30; // @[HandShaking.scala 232:72]
  wire  _T_31; // @[HandShaking.scala 232:72]
  wire  _T_32; // @[ComputeNode.scala 107:17]
  wire  _T_33; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_23_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_18; // @[ComputeNode.scala 99:61]
  wire  _GEN_27; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _GEN_29; // @[ComputeNode.scala 99:61]
  wire  _GEN_35; // @[ComputeNode.scala 99:61]
  wire  _T_38; // @[HandShaking.scala 217:83]
  wire  _T_39; // @[HandShaking.scala 217:83]
  wire  _T_40; // @[HandShaking.scala 217:83]
  wire  _T_41; // @[HandShaking.scala 218:27]
  wire  _T_42; // @[HandShaking.scala 218:27]
  wire  _GEN_71; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _T_5 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_14 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_16 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_16 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_20 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_22 = _T_21 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_29 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_30 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_31 = _T_3 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_32 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_33 = _T_32 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_23_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_18 = _T_22 ? _T_23_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_27 = _T_22 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_22 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_29 = _T_22 | out_valid_R_2; // @[ComputeNode.scala 99:61]
  assign _GEN_35 = _T_22 | state; // @[ComputeNode.scala 99:61]
  assign _T_38 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_39 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_40 = out_ready_R_2 | _T_3; // @[HandShaking.scala 217:83]
  assign _T_41 = _T_38 & _T_39; // @[HandShaking.scala 218:27]
  assign _T_42 = _T_41 & _T_40; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_20 ? _GEN_27 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_20 ? _GEN_18 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_20 ? _GEN_28 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_20 ? _GEN_18 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_2_valid = _T_20 ? _GEN_29 : out_valid_R_2; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_2_bits_data = _T_20 ? _GEN_18 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_71 = _T_20 & _T_22; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value = _RAND_9[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  left_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  left_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  right_R_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  right_valid_R = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_data_R = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_5) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_5) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_5) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_5) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_5) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_3) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          out_valid_R_0 <= _T_29;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          out_valid_R_1 <= _T_30;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          out_valid_R_2 <= _T_31;
        end else begin
          if (_T_3) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_3) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_8;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_13;
        end
      end else begin
        left_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_16) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_17;
        end
      end else begin
        right_valid_R <= _GEN_17;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_20) begin
        state <= _GEN_35;
      end else begin
        if (state) begin
          if (_T_42) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_20) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & _T_33) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add5358: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_12(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx5459: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_8(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_60: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_60: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_60: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ZextNode_3(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[ZextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[ZextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[ZextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[ZextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[ZextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[ZextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[ZextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[ZextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[ZextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[ZextNode.scala 84:26]
  wire  _GEN_9; // @[ZextNode.scala 84:26]
  wire  fire_mask_0; // @[ZextNode.scala 90:74]
  reg  state; // @[ZextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[ZextNode.scala 93:27]
  wire  _T_16; // @[ZextNode.scala 97:26]
  wire  _T_17; // @[ZextNode.scala 110:28]
  wire  _T_18; // @[ZextNode.scala 117:17]
  wire  _T_19; // @[ZextNode.scala 117:17]
  wire  _GEN_10; // @[ZextNode.scala 110:47]
  wire  _GEN_11; // @[ZextNode.scala 110:47]
  wire  _GEN_42; // @[ZextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ZextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[ZextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[ZextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[ZextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[ZextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[ZextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[ZextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[ZextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[ZextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[ZextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[ZextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[ZextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[ZextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[ZextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[ZextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[ZextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[ZextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[ZextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] sextconv5661: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[ZextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_27(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul5762: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_28(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add5863: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore_3(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [STORE]st_64: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_9(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_65: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_65: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_65: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_29(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add6566: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_13(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx6667: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_10(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_68: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_68: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_68: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ZextNode_4(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[ZextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[ZextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[ZextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[ZextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[ZextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[ZextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[ZextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[ZextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[ZextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[ZextNode.scala 84:26]
  wire  _GEN_9; // @[ZextNode.scala 84:26]
  wire  fire_mask_0; // @[ZextNode.scala 90:74]
  reg  state; // @[ZextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[ZextNode.scala 93:27]
  wire  _T_16; // @[ZextNode.scala 97:26]
  wire  _T_17; // @[ZextNode.scala 110:28]
  wire  _T_18; // @[ZextNode.scala 117:17]
  wire  _T_19; // @[ZextNode.scala 117:17]
  wire  _GEN_10; // @[ZextNode.scala 110:47]
  wire  _GEN_11; // @[ZextNode.scala 110:47]
  wire  _GEN_42; // @[ZextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ZextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[ZextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[ZextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[ZextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[ZextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[ZextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[ZextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[ZextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[ZextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[ZextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[ZextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[ZextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[ZextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[ZextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[ZextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[ZextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[ZextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[ZextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] sextconv6869: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[ZextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_30(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul6970: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_31(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add7071: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore_4(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [STORE]st_72: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_11(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_73: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_73: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_73: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_32(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h2;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add7774: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_14(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx7875: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_12(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_76: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_76: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_76: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ZextNode_5(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[ZextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[ZextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[ZextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[ZextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[ZextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[ZextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[ZextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[ZextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[ZextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[ZextNode.scala 84:26]
  wire  _GEN_9; // @[ZextNode.scala 84:26]
  wire  fire_mask_0; // @[ZextNode.scala 90:74]
  reg  state; // @[ZextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[ZextNode.scala 93:27]
  wire  _T_16; // @[ZextNode.scala 97:26]
  wire  _T_17; // @[ZextNode.scala 110:28]
  wire  _T_18; // @[ZextNode.scala 117:17]
  wire  _T_19; // @[ZextNode.scala 117:17]
  wire  _GEN_10; // @[ZextNode.scala 110:47]
  wire  _GEN_11; // @[ZextNode.scala 110:47]
  wire  _GEN_42; // @[ZextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ZextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[ZextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[ZextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[ZextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[ZextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[ZextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[ZextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[ZextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[ZextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[ZextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[ZextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[ZextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[ZextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[ZextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[ZextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[ZextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[ZextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[ZextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] sextconv8077: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[ZextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_33(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul8178: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_34(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add8279: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore_5(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [STORE]st_80: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_13(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_81: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_81: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_81: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_35(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  input         io_Out_2_ready,
  output        io_Out_2_valid,
  output [31:0] io_Out_2_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_ready_R_2; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_7;
  reg  out_valid_R_2; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_8;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  wire  _T_5; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_9;
  wire [14:0] _T_8; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_10;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_11;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_12;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_13;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_14;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_15;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 74:26]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_17; // @[ComputeNode.scala 80:27]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[ComputeNode.scala 99:27]
  wire  _T_22; // @[ComputeNode.scala 99:43]
  wire  _T_29; // @[HandShaking.scala 232:72]
  wire  _T_30; // @[HandShaking.scala 232:72]
  wire  _T_31; // @[HandShaking.scala 232:72]
  wire  _T_32; // @[ComputeNode.scala 107:17]
  wire  _T_33; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_23_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_18; // @[ComputeNode.scala 99:61]
  wire  _GEN_27; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _GEN_29; // @[ComputeNode.scala 99:61]
  wire  _GEN_35; // @[ComputeNode.scala 99:61]
  wire  _T_38; // @[HandShaking.scala 217:83]
  wire  _T_39; // @[HandShaking.scala 217:83]
  wire  _T_40; // @[HandShaking.scala 217:83]
  wire  _T_41; // @[HandShaking.scala 218:27]
  wire  _T_42; // @[HandShaking.scala 218:27]
  wire  _GEN_71; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_Out_2_ready & io_Out_2_valid; // @[Decoupled.scala 40:37]
  assign _T_5 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_8 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_14 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_16 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_17 = _T_16 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_20 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_22 = _T_21 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_29 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_30 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_31 = _T_3 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_32 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_33 = _T_32 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_23_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_18 = _T_22 ? _T_23_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_27 = _T_22 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_22 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_29 = _T_22 | out_valid_R_2; // @[ComputeNode.scala 99:61]
  assign _GEN_35 = _T_22 | state; // @[ComputeNode.scala 99:61]
  assign _T_38 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_39 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_40 = out_ready_R_2 | _T_3; // @[HandShaking.scala 217:83]
  assign _T_41 = _T_38 & _T_39; // @[HandShaking.scala 218:27]
  assign _T_42 = _T_41 & _T_40; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_20 ? _GEN_27 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_20 ? _GEN_18 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_20 ? _GEN_28 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_20 ? _GEN_18 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_2_valid = _T_20 ? _GEN_29 : out_valid_R_2; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_2_bits_data = _T_20 ? _GEN_18 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_71 = _T_20 & _T_22; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_ready_R_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  out_valid_R_2 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  value = _RAND_9[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  left_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  left_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  right_R_data = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  right_valid_R = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  out_data_R = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_5) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_5) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_5) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_5) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_5) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_2 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_3) begin
          out_ready_R_2 <= io_Out_2_ready;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_ready_R_2 <= 1'h0;
          end else begin
            if (_T_3) begin
              out_ready_R_2 <= io_Out_2_ready;
            end
          end
        end else begin
          if (_T_3) begin
            out_ready_R_2 <= io_Out_2_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          out_valid_R_0 <= _T_29;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          out_valid_R_1 <= _T_30;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_2 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          out_valid_R_2 <= _T_31;
        end else begin
          if (_T_3) begin
            out_valid_R_2 <= 1'h0;
          end
        end
      end else begin
        if (_T_3) begin
          out_valid_R_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_8;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_13;
        end
      end else begin
        left_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_16) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_22) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_17;
        end
      end else begin
        right_valid_R <= _GEN_17;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_20) begin
        state <= _GEN_35;
      end else begin
        if (state) begin
          if (_T_42) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_20) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_42) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_71 & _T_33) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add8882: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_15(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx8983: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_14(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_84: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_84: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_84: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ZextNode_6(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[ZextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[ZextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[ZextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[ZextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[ZextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[ZextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[ZextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[ZextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[ZextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[ZextNode.scala 84:26]
  wire  _GEN_9; // @[ZextNode.scala 84:26]
  wire  fire_mask_0; // @[ZextNode.scala 90:74]
  reg  state; // @[ZextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[ZextNode.scala 93:27]
  wire  _T_16; // @[ZextNode.scala 97:26]
  wire  _T_17; // @[ZextNode.scala 110:28]
  wire  _T_18; // @[ZextNode.scala 117:17]
  wire  _T_19; // @[ZextNode.scala 117:17]
  wire  _GEN_10; // @[ZextNode.scala 110:47]
  wire  _GEN_11; // @[ZextNode.scala 110:47]
  wire  _GEN_42; // @[ZextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ZextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[ZextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[ZextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[ZextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[ZextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[ZextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[ZextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[ZextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[ZextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[ZextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[ZextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[ZextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[ZextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[ZextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[ZextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[ZextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[ZextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[ZextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] sextconv9185: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[ZextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_36(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul9286: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_37(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add9387: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore_6(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [STORE]st_88: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_15(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_89: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_89: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_89: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_38(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add10090: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_16(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx10191: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_16(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_92: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_92: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_92: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ZextNode_7(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[ZextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[ZextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[ZextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[ZextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[ZextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[ZextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[ZextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[ZextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[ZextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[ZextNode.scala 84:26]
  wire  _GEN_9; // @[ZextNode.scala 84:26]
  wire  fire_mask_0; // @[ZextNode.scala 90:74]
  reg  state; // @[ZextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[ZextNode.scala 93:27]
  wire  _T_16; // @[ZextNode.scala 97:26]
  wire  _T_17; // @[ZextNode.scala 110:28]
  wire  _T_18; // @[ZextNode.scala 117:17]
  wire  _T_19; // @[ZextNode.scala 117:17]
  wire  _GEN_10; // @[ZextNode.scala 110:47]
  wire  _GEN_11; // @[ZextNode.scala 110:47]
  wire  _GEN_42; // @[ZextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ZextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[ZextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[ZextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[ZextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[ZextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[ZextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[ZextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[ZextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[ZextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[ZextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[ZextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[ZextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[ZextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[ZextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[ZextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[ZextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[ZextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[ZextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] sextconv10393: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[ZextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_39(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul10494: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_40(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add10595: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore_7(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [STORE]st_96: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_17(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_97: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_97: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_97: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_41(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h2;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add11298: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module GepNode_17(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output        io_Out_0_bits_predicate,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_baseAddress_ready,
  input         io_baseAddress_valid,
  input  [4:0]  io_baseAddress_bits_taskID,
  input  [31:0] io_baseAddress_bits_data,
  output        io_idx_0_ready,
  input         io_idx_0_valid,
  input  [31:0] io_idx_0_bits_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [4:0] base_addr_R_taskID; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_6;
  reg [31:0] base_addr_R_data; // @[GepNode.scala 880:28]
  reg [31:0] _RAND_7;
  reg  base_addr_valid_R; // @[GepNode.scala 881:34]
  reg [31:0] _RAND_8;
  reg [31:0] idx_R_0_data; // @[GepNode.scala 884:39]
  reg [31:0] _RAND_9;
  reg  idx_valid_R_0; // @[GepNode.scala 885:45]
  reg [31:0] _RAND_10;
  reg  state; // @[GepNode.scala 889:22]
  reg [31:0] _RAND_11;
  wire  _T_11; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[GepNode.scala 905:31]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[GepNode.scala 912:28]
  wire [32:0] seek_value; // @[GepNode.scala 920:21]
  wire [32:0] _GEN_50; // @[GepNode.scala 928:35]
  wire [32:0] data_out; // @[GepNode.scala 928:35]
  wire  _T_15; // @[Conditional.scala 37:30]
  wire  _T_16; // @[GepNode.scala 944:27]
  wire  _T_17; // @[GepNode.scala 944:48]
  wire  _T_19; // @[HandShaking.scala 232:72]
  wire  _GEN_15; // @[GepNode.scala 944:78]
  wire  _T_22; // @[HandShaking.scala 217:83]
  wire  _T_25; // @[GepNode.scala 964:17]
  wire  _T_26; // @[GepNode.scala 964:17]
  wire  _GEN_51; // @[GepNode.scala 964:17]
  wire  _GEN_52; // @[GepNode.scala 964:17]
  wire  _GEN_53; // @[GepNode.scala 964:17]
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_11 = io_baseAddress_ready & io_baseAddress_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_11 | base_addr_valid_R; // @[GepNode.scala 905:31]
  assign _T_13 = io_idx_0_ready & io_idx_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_13 | idx_valid_R_0; // @[GepNode.scala 912:28]
  assign seek_value = idx_R_0_data * 32'h1; // @[GepNode.scala 920:21]
  assign _GEN_50 = {{1'd0}, base_addr_R_data}; // @[GepNode.scala 928:35]
  assign data_out = _GEN_50 + seek_value; // @[GepNode.scala 928:35]
  assign _T_15 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_16 = enable_valid_R & base_addr_valid_R; // @[GepNode.scala 944:27]
  assign _T_17 = _T_16 & idx_valid_R_0; // @[GepNode.scala 944:48]
  assign _T_19 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _GEN_15 = _T_17 | state; // @[GepNode.scala 944:78]
  assign _T_22 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_25 = $unsigned(reset); // @[GepNode.scala 964:17]
  assign _T_26 = _T_25 == 1'h0; // @[GepNode.scala 964:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 180:21]
  assign io_Out_0_bits_predicate = enable_R_control; // @[GepNode.scala 933:30]
  assign io_Out_0_bits_taskID = base_addr_R_taskID; // @[GepNode.scala 934:27]
  assign io_Out_0_bits_data = data_out[31:0]; // @[GepNode.scala 932:25]
  assign io_baseAddress_ready = ~ base_addr_valid_R; // @[GepNode.scala 904:24]
  assign io_idx_0_ready = ~ idx_valid_R_0; // @[GepNode.scala 911:21]
  assign _GEN_51 = _T_15 == 1'h0; // @[GepNode.scala 964:17]
  assign _GEN_52 = _GEN_51 & state; // @[GepNode.scala 964:17]
  assign _GEN_53 = _GEN_52 & _T_22; // @[GepNode.scala 964:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  base_addr_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  base_addr_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  base_addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  idx_R_0_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  idx_valid_R_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        if (_T_17) begin
          out_valid_R_0 <= _T_19;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      base_addr_R_taskID <= 5'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_taskID <= io_baseAddress_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_taskID <= 5'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_taskID <= io_baseAddress_bits_taskID;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_taskID <= io_baseAddress_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      base_addr_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_11) begin
          base_addr_R_data <= io_baseAddress_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_R_data <= 32'h0;
          end else begin
            if (_T_11) begin
              base_addr_R_data <= io_baseAddress_bits_data;
            end
          end
        end else begin
          if (_T_11) begin
            base_addr_R_data <= io_baseAddress_bits_data;
          end
        end
      end
    end
    if (reset) begin
      base_addr_valid_R <= 1'h0;
    end else begin
      if (_T_15) begin
        base_addr_valid_R <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_22) begin
            base_addr_valid_R <= 1'h0;
          end else begin
            base_addr_valid_R <= _GEN_9;
          end
        end else begin
          base_addr_valid_R <= _GEN_9;
        end
      end
    end
    if (reset) begin
      idx_R_0_data <= 32'h0;
    end else begin
      if (_T_15) begin
        if (_T_13) begin
          idx_R_0_data <= io_idx_0_bits_data;
        end
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_R_0_data <= 32'h0;
          end else begin
            if (_T_13) begin
              idx_R_0_data <= io_idx_0_bits_data;
            end
          end
        end else begin
          if (_T_13) begin
            idx_R_0_data <= io_idx_0_bits_data;
          end
        end
      end
    end
    if (reset) begin
      idx_valid_R_0 <= 1'h0;
    end else begin
      if (_T_15) begin
        idx_valid_R_0 <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_22) begin
            idx_valid_R_0 <= 1'h0;
          end else begin
            idx_valid_R_0 <= _GEN_13;
          end
        end else begin
          idx_valid_R_0 <= _GEN_13;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_15) begin
        state <= _GEN_15;
      end else begin
        if (state) begin
          if (_T_22) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_53 & _T_26) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [GEP] Gep_arrayidx11399: Output fired @ %d, Value: %d\n",enable_R_taskID,value,data_out); // @[GepNode.scala 964:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypLoad_18(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input         io_GepAddr_bits_predicate,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [31:0] io_memReq_bits_address,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid,
  input  [31:0] io_memResp_data
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 530:28]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 531:28]
  reg [31:0] _RAND_4;
  wire  _T_4; // @[Decoupled.scala 40:37]
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg  addr_R_predicate; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_6;
  reg [4:0] addr_R_taskID; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_7;
  reg [31:0] addr_R_data; // @[LoadSimple.scala 63:23]
  reg [31:0] _RAND_8;
  reg  addr_valid_R; // @[LoadSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [31:0] data_R_data; // @[LoadSimple.scala 67:23]
  reg [31:0] _RAND_10;
  reg [1:0] state; // @[LoadSimple.scala 72:22]
  reg [31:0] _RAND_11;
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[LoadSimple.scala 81:27]
  wire  complete; // @[HandShaking.scala 648:29]
  wire  predicate; // @[LoadSimple.scala 91:36]
  wire  _T_20; // @[Conditional.scala 37:30]
  wire  _T_21; // @[LoadSimple.scala 119:27]
  wire  _T_22; // @[LoadSimple.scala 120:31]
  wire  _T_23; // @[Decoupled.scala 40:37]
  wire  _T_24; // @[LoadSimple.scala 125:21]
  wire  _T_25; // @[LoadSimple.scala 125:21]
  wire  _T_27; // @[HandShaking.scala 652:72]
  wire  _GEN_15; // @[LoadSimple.scala 119:44]
  wire  _T_28; // @[Conditional.scala 37:30]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _GEN_50; // @[LoadSimple.scala 125:21]
  wire  _GEN_51; // @[LoadSimple.scala 125:21]
  wire  _GEN_52; // @[LoadSimple.scala 125:21]
  wire  _GEN_53; // @[LoadSimple.scala 151:17]
  wire  _GEN_54; // @[LoadSimple.scala 151:17]
  wire  _GEN_55; // @[LoadSimple.scala 151:17]
  wire  _GEN_57; // @[LoadSimple.scala 172:17]
  wire  _GEN_58; // @[LoadSimple.scala 172:17]
  wire  _GEN_59; // @[LoadSimple.scala 172:17]
  wire  _GEN_60; // @[LoadSimple.scala 172:17]
  assign _T_4 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_14 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_14 | addr_valid_R; // @[LoadSimple.scala 81:27]
  assign complete = out_ready_R_0 | io_Out_0_ready; // @[HandShaking.scala 648:29]
  assign predicate = addr_R_predicate & enable_R_control; // @[LoadSimple.scala 91:36]
  assign _T_20 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_21 = enable_valid_R & addr_valid_R; // @[LoadSimple.scala 119:27]
  assign _T_22 = enable_R_control & predicate; // @[LoadSimple.scala 120:31]
  assign _T_23 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _T_24 = $unsigned(reset); // @[LoadSimple.scala 125:21]
  assign _T_25 = _T_24 == 1'h0; // @[LoadSimple.scala 125:21]
  assign _T_27 = _T_4 ^ 1'h1; // @[HandShaking.scala 652:72]
  assign _GEN_15 = _T_21 & _T_22; // @[LoadSimple.scala 119:44]
  assign _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_Out_0_valid = out_valid_R_0; // @[HandShaking.scala 555:21]
  assign io_Out_0_bits_data = data_R_data; // @[LoadSimple.scala 97:20]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[LoadSimple.scala 80:20]
  assign io_memReq_valid = _T_20 & _GEN_15; // @[LoadSimple.scala 102:19 LoadSimple.scala 121:27]
  assign io_memReq_bits_address = addr_R_data; // @[LoadSimple.scala 103:26]
  assign io_memReq_bits_taskID = addr_R_taskID; // @[LoadSimple.scala 106:25]
  assign _GEN_50 = _T_20 & _T_21; // @[LoadSimple.scala 125:21]
  assign _GEN_51 = _GEN_50 & _T_22; // @[LoadSimple.scala 125:21]
  assign _GEN_52 = _GEN_51 & _T_23; // @[LoadSimple.scala 125:21]
  assign _GEN_53 = _T_20 == 1'h0; // @[LoadSimple.scala 151:17]
  assign _GEN_54 = _GEN_53 & _T_28; // @[LoadSimple.scala 151:17]
  assign _GEN_55 = _GEN_54 & io_memResp_valid; // @[LoadSimple.scala 151:17]
  assign _GEN_57 = _T_28 == 1'h0; // @[LoadSimple.scala 172:17]
  assign _GEN_58 = _GEN_53 & _GEN_57; // @[LoadSimple.scala 172:17]
  assign _GEN_59 = _GEN_58 & _T_33; // @[LoadSimple.scala 172:17]
  assign _GEN_60 = _GEN_59 & complete; // @[LoadSimple.scala 172:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  addr_R_predicate = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  addr_R_taskID = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  addr_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  data_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  state = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_28) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              enable_valid_R <= 1'h0;
            end else begin
              if (_T_6) begin
                enable_valid_R <= io_enable_valid;
              end
            end
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_4) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (_T_28) begin
          if (_T_4) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              out_ready_R_0 <= 1'h0;
            end else begin
              if (_T_4) begin
                out_ready_R_0 <= io_Out_0_ready;
              end
            end
          end else begin
            if (_T_4) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end else begin
            out_valid_R_0 <= _T_27;
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            out_valid_R_0 <= _T_27;
          end else begin
            if (_T_4) begin
              out_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_4) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_predicate <= 1'h0;
    end else begin
      if (_T_14) begin
        addr_R_predicate <= io_GepAddr_bits_predicate;
      end
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_14) begin
        addr_R_taskID <= io_GepAddr_bits_taskID;
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        addr_R_data <= io_GepAddr_bits_data;
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_20) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_28) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_33) begin
            if (complete) begin
              addr_valid_R <= 1'h0;
            end else begin
              addr_valid_R <= _GEN_9;
            end
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (!(_T_20)) begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            data_R_data <= io_memResp_data;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_20) begin
        if (_T_21) begin
          if (_T_22) begin
            if (_T_23) begin
              state <= 2'h1;
            end
          end else begin
            state <= 2'h2;
          end
        end
      end else begin
        if (_T_28) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_33) begin
            if (complete) begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_52 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_100: Memreq fired @ %d, Addr:%d\n",enable_R_taskID,value,io_memReq_bits_address); // @[LoadSimple.scala 125:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_55 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_100: Memresp fired @ %d, Value: %d\n",enable_R_taskID,value,io_memResp_data); // @[LoadSimple.scala 151:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_25) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [LOAD] ld_100: Output fired @ %d, Address:%d, Value: %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[LoadSimple.scala 172:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ZextNode_8(
  input         clock,
  input         reset,
  output        io_Input_ready,
  input         io_Input_valid,
  input  [31:0] io_Input_bits_data,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [31:0] input_R_data; // @[ZextNode.scala 47:24]
  reg [31:0] _RAND_1;
  reg  input_valid_R; // @[ZextNode.scala 48:30]
  reg [31:0] _RAND_2;
  reg [4:0] enable_R_taskID; // @[ZextNode.scala 50:25]
  reg [31:0] _RAND_3;
  reg  enable_valid_R; // @[ZextNode.scala 51:31]
  reg [31:0] _RAND_4;
  reg  output_valid_R_0; // @[ZextNode.scala 53:49]
  reg [31:0] _RAND_5;
  reg  fire_R_0; // @[ZextNode.scala 55:41]
  reg [31:0] _RAND_6;
  wire [4:0] task_input; // @[ZextNode.scala 57:43]
  wire  _T_7; // @[Decoupled.scala 40:37]
  wire  _GEN_4; // @[ZextNode.scala 65:25]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[ZextNode.scala 71:26]
  wire  _T_10; // @[Decoupled.scala 40:37]
  wire  _GEN_8; // @[ZextNode.scala 84:26]
  wire  _GEN_9; // @[ZextNode.scala 84:26]
  wire  fire_mask_0; // @[ZextNode.scala 90:74]
  reg  state; // @[ZextNode.scala 105:22]
  reg [31:0] _RAND_7;
  wire  _T_12; // @[Conditional.scala 37:30]
  wire  _T_14; // @[ZextNode.scala 93:27]
  wire  _T_16; // @[ZextNode.scala 97:26]
  wire  _T_17; // @[ZextNode.scala 110:28]
  wire  _T_18; // @[ZextNode.scala 117:17]
  wire  _T_19; // @[ZextNode.scala 117:17]
  wire  _GEN_10; // @[ZextNode.scala 110:47]
  wire  _GEN_11; // @[ZextNode.scala 110:47]
  wire  _GEN_42; // @[ZextNode.scala 117:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_input = io_enable_bits_taskID | enable_R_taskID; // @[ZextNode.scala 57:43]
  assign _T_7 = io_Input_ready & io_Input_valid; // @[Decoupled.scala 40:37]
  assign _GEN_4 = _T_7 | input_valid_R; // @[ZextNode.scala 65:25]
  assign _T_9 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_9 | enable_valid_R; // @[ZextNode.scala 71:26]
  assign _T_10 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_8 = _T_10 ? 1'h0 : output_valid_R_0; // @[ZextNode.scala 84:26]
  assign _GEN_9 = _T_10 | fire_R_0; // @[ZextNode.scala 84:26]
  assign fire_mask_0 = fire_R_0 | _T_10; // @[ZextNode.scala 90:74]
  assign _T_12 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_14 = enable_valid_R | _T_9; // @[ZextNode.scala 93:27]
  assign _T_16 = input_valid_R | _T_7; // @[ZextNode.scala 97:26]
  assign _T_17 = _T_14 & _T_16; // @[ZextNode.scala 110:28]
  assign _T_18 = $unsigned(reset); // @[ZextNode.scala 117:17]
  assign _T_19 = _T_18 == 1'h0; // @[ZextNode.scala 117:17]
  assign _GEN_10 = _T_17 | _GEN_8; // @[ZextNode.scala 110:47]
  assign _GEN_11 = _T_17 | state; // @[ZextNode.scala 110:47]
  assign io_Input_ready = ~ input_valid_R; // @[ZextNode.scala 64:18]
  assign io_enable_ready = ~ enable_valid_R; // @[ZextNode.scala 70:19]
  assign io_Out_0_valid = output_valid_R_0; // @[ZextNode.scala 80:21]
  assign io_Out_0_bits_data = input_R_data; // @[ZextNode.scala 79:20]
  assign _GEN_42 = _T_12 & _T_17; // @[ZextNode.scala 117:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  input_R_data = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  input_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  enable_R_taskID = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_valid_R = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  output_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  fire_R_0 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  state = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      input_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        if (_T_7) begin
          input_R_data <= io_Input_bits_data;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_R_data <= 32'h0;
          end else begin
            if (_T_7) begin
              input_R_data <= io_Input_bits_data;
            end
          end
        end else begin
          if (_T_7) begin
            input_R_data <= io_Input_bits_data;
          end
        end
      end
    end
    if (reset) begin
      input_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        input_valid_R <= _GEN_4;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            input_valid_R <= 1'h0;
          end else begin
            input_valid_R <= _GEN_4;
          end
        end else begin
          input_valid_R <= _GEN_4;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_12) begin
        if (_T_9) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_12) begin
        enable_valid_R <= _GEN_7;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_7;
          end
        end else begin
          enable_valid_R <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_valid_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        output_valid_R_0 <= _GEN_10;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            output_valid_R_0 <= 1'h0;
          end else begin
            if (_T_10) begin
              output_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_10) begin
            output_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_R_0 <= 1'h0;
    end else begin
      if (_T_12) begin
        fire_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            fire_R_0 <= 1'h0;
          end else begin
            fire_R_0 <= _GEN_9;
          end
        end else begin
          fire_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_12) begin
        state <= _GEN_11;
      end else begin
        if (state) begin
          if (fire_mask_0) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_42 & _T_19) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] sextconv115101: Output fired @ %d, Value: %d\n",task_input,value,input_R_data); // @[ZextNode.scala 117:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_42(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_mul116102: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_43(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid,
  input  [31:0] io_RightIO_bits_data
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= io_RightIO_bits_data;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_add117103: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module UnTypStore_8(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_GepAddr_ready,
  input         io_GepAddr_valid,
  input  [4:0]  io_GepAddr_bits_taskID,
  input  [31:0] io_GepAddr_bits_data,
  output        io_inData_ready,
  input         io_inData_valid,
  input  [4:0]  io_inData_bits_taskID,
  input  [31:0] io_inData_bits_data,
  input         io_memReq_ready,
  output        io_memReq_valid,
  output [21:0] io_memReq_bits_address,
  output [31:0] io_memReq_bits_data,
  output [4:0]  io_memReq_bits_taskID,
  input         io_memResp_valid
);
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 517:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 518:31]
  reg [31:0] _RAND_2;
  wire  _T_6; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_3;
  wire [14:0] _T_9; // @[Counter.scala 38:22]
  reg [4:0] addr_R_taskID; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_4;
  reg [31:0] addr_R_data; // @[StoreSimple.scala 61:23]
  reg [31:0] _RAND_5;
  reg [4:0] data_R_taskID; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_6;
  reg [31:0] data_R_data; // @[StoreSimple.scala 62:23]
  reg [31:0] _RAND_7;
  reg  addr_valid_R; // @[StoreSimple.scala 63:29]
  reg [31:0] _RAND_8;
  reg  data_valid_R; // @[StoreSimple.scala 64:29]
  reg [31:0] _RAND_9;
  reg [1:0] state; // @[StoreSimple.scala 68:22]
  reg [31:0] _RAND_10;
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[StoreSimple.scala 89:27]
  wire  _T_18; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[StoreSimple.scala 97:26]
  wire [4:0] _T_19; // @[StoreSimple.scala 106:44]
  wire  mem_req_fire; // @[StoreSimple.scala 120:51]
  wire  _T_27; // @[Conditional.scala 37:30]
  wire  _T_28; // @[StoreSimple.scala 126:27]
  wire  _T_29; // @[StoreSimple.scala 127:33]
  wire  _T_30; // @[Decoupled.scala 40:37]
  wire  _GEN_19; // @[StoreSimple.scala 126:44]
  wire  _GEN_23; // @[StoreSimple.scala 125:28]
  wire  _T_33; // @[Conditional.scala 37:30]
  wire  _T_36; // @[Conditional.scala 37:30]
  wire  _T_40; // @[StoreSimple.scala 162:17]
  wire  _T_41; // @[StoreSimple.scala 162:17]
  wire  _GEN_76; // @[StoreSimple.scala 162:17]
  wire  _GEN_77; // @[StoreSimple.scala 162:17]
  wire  _GEN_78; // @[StoreSimple.scala 162:17]
  wire  _GEN_79; // @[StoreSimple.scala 162:17]
  assign _T_6 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = value + 15'h1; // @[Counter.scala 38:22]
  assign _T_16 = io_GepAddr_ready & io_GepAddr_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | addr_valid_R; // @[StoreSimple.scala 89:27]
  assign _T_18 = io_inData_ready & io_inData_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_18 | data_valid_R; // @[StoreSimple.scala 97:26]
  assign _T_19 = data_R_taskID | addr_R_taskID; // @[StoreSimple.scala 106:44]
  assign mem_req_fire = addr_valid_R & data_valid_R; // @[StoreSimple.scala 120:51]
  assign _T_27 = 2'h0 == state; // @[Conditional.scala 37:30]
  assign _T_28 = data_valid_R & addr_valid_R; // @[StoreSimple.scala 126:27]
  assign _T_29 = enable_R_control & mem_req_fire; // @[StoreSimple.scala 127:33]
  assign _T_30 = io_memReq_ready & io_memReq_valid; // @[Decoupled.scala 40:37]
  assign _GEN_19 = _T_28 & _T_29; // @[StoreSimple.scala 126:44]
  assign _GEN_23 = enable_valid_R & _GEN_19; // @[StoreSimple.scala 125:28]
  assign _T_33 = 2'h1 == state; // @[Conditional.scala 37:30]
  assign _T_36 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign _T_40 = $unsigned(reset); // @[StoreSimple.scala 162:17]
  assign _T_41 = _T_40 == 1'h0; // @[StoreSimple.scala 162:17]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 575:19]
  assign io_GepAddr_ready = ~ addr_valid_R; // @[StoreSimple.scala 84:20 StoreSimple.scala 88:20]
  assign io_inData_ready = ~ data_valid_R; // @[StoreSimple.scala 85:19]
  assign io_memReq_valid = _T_27 & _GEN_23; // @[StoreSimple.scala 115:19 StoreSimple.scala 128:29]
  assign io_memReq_bits_address = addr_R_data[21:0]; // @[StoreSimple.scala 109:26]
  assign io_memReq_bits_data = data_R_data; // @[StoreSimple.scala 110:23]
  assign io_memReq_bits_taskID = _T_19 | enable_R_taskID; // @[StoreSimple.scala 113:25]
  assign _GEN_76 = _T_27 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_77 = _T_33 == 1'h0; // @[StoreSimple.scala 162:17]
  assign _GEN_78 = _GEN_76 & _GEN_77; // @[StoreSimple.scala 162:17]
  assign _GEN_79 = _GEN_78 & _T_36; // @[StoreSimple.scala 162:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  addr_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  addr_R_data = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  data_R_taskID = _RAND_6[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  data_R_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr_valid_R = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  data_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_6) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_6) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        if (_T_6) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (_T_33) begin
          if (_T_6) begin
            enable_valid_R <= io_enable_valid;
          end
        end else begin
          if (_T_36) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_6) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_9;
    end
    if (reset) begin
      addr_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_taskID <= io_GepAddr_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_taskID <= io_GepAddr_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            addr_R_taskID <= 5'h0;
          end else begin
            if (_T_16) begin
              addr_R_taskID <= io_GepAddr_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_16) begin
          addr_R_data <= io_GepAddr_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_16) begin
            addr_R_data <= io_GepAddr_bits_data;
          end
        end else begin
          if (_T_36) begin
            addr_R_data <= 32'h0;
          end else begin
            if (_T_16) begin
              addr_R_data <= io_GepAddr_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_taskID <= 5'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_taskID <= io_inData_bits_taskID;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_taskID <= io_inData_bits_taskID;
          end
        end else begin
          if (_T_36) begin
            data_R_taskID <= 5'h0;
          end else begin
            if (_T_18) begin
              data_R_taskID <= io_inData_bits_taskID;
            end
          end
        end
      end
    end
    if (reset) begin
      data_R_data <= 32'h0;
    end else begin
      if (_T_27) begin
        if (_T_18) begin
          data_R_data <= io_inData_bits_data;
        end
      end else begin
        if (_T_33) begin
          if (_T_18) begin
            data_R_data <= io_inData_bits_data;
          end
        end else begin
          if (_T_36) begin
            data_R_data <= 32'h0;
          end else begin
            if (_T_18) begin
              data_R_data <= io_inData_bits_data;
            end
          end
        end
      end
    end
    if (reset) begin
      addr_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        addr_valid_R <= _GEN_9;
      end else begin
        if (_T_33) begin
          addr_valid_R <= _GEN_9;
        end else begin
          if (_T_36) begin
            addr_valid_R <= 1'h0;
          end else begin
            addr_valid_R <= _GEN_9;
          end
        end
      end
    end
    if (reset) begin
      data_valid_R <= 1'h0;
    end else begin
      if (_T_27) begin
        data_valid_R <= _GEN_13;
      end else begin
        if (_T_33) begin
          data_valid_R <= _GEN_13;
        end else begin
          if (_T_36) begin
            data_valid_R <= 1'h0;
          end else begin
            data_valid_R <= _GEN_13;
          end
        end
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_27) begin
        if (enable_valid_R) begin
          if (_T_28) begin
            if (_T_29) begin
              if (_T_30) begin
                state <= 2'h1;
              end
            end else begin
              state <= 2'h2;
            end
          end
        end
      end else begin
        if (_T_33) begin
          if (io_memResp_valid) begin
            state <= 2'h2;
          end
        end else begin
          if (_T_36) begin
            state <= 2'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_79 & _T_41) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [STORE]st_104: Fired @ %d Mem[%d] = %d\n",enable_R_taskID,value,addr_R_data,data_R_data); // @[StoreSimple.scala 162:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_44(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  input         io_Out_1_ready,
  output        io_Out_1_valid,
  output [31:0] io_Out_1_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_ready_R_1; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_4;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_5;
  reg  out_valid_R_1; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_6;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_2; // @[Decoupled.scala 40:37]
  wire  _T_4; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_7;
  wire [14:0] _T_7; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_8;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_9;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_10;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_11;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_12;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_13;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_13; // @[Decoupled.scala 40:37]
  wire  _GEN_11; // @[ComputeNode.scala 74:26]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_15; // @[ComputeNode.scala 80:27]
  wire  _T_18; // @[Conditional.scala 37:30]
  wire  _T_19; // @[ComputeNode.scala 99:27]
  wire  _T_20; // @[ComputeNode.scala 99:43]
  wire  _T_25; // @[HandShaking.scala 232:72]
  wire  _T_26; // @[HandShaking.scala 232:72]
  wire  _T_27; // @[ComputeNode.scala 107:17]
  wire  _T_28; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_21_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_16; // @[ComputeNode.scala 99:61]
  wire  _GEN_22; // @[ComputeNode.scala 99:61]
  wire  _GEN_23; // @[ComputeNode.scala 99:61]
  wire  _GEN_28; // @[ComputeNode.scala 99:61]
  wire  _T_32; // @[HandShaking.scala 217:83]
  wire  _T_33; // @[HandShaking.scala 217:83]
  wire  _T_34; // @[HandShaking.scala 218:27]
  wire  _GEN_56; // @[ComputeNode.scala 107:17]
  UALU_1 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_2 = io_Out_1_ready & io_Out_1_valid; // @[Decoupled.scala 40:37]
  assign _T_4 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_7 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_13 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_11 = _T_13 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_15 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_15 = _T_15 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_18 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_19 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_20 = _T_19 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_25 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_26 = _T_2 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_27 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_28 = _T_27 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_21_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_16 = _T_20 ? _T_21_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_22 = _T_20 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_23 = _T_20 | out_valid_R_1; // @[ComputeNode.scala 99:61]
  assign _GEN_28 = _T_20 | state; // @[ComputeNode.scala 99:61]
  assign _T_32 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign _T_33 = out_ready_R_1 | _T_2; // @[HandShaking.scala 217:83]
  assign _T_34 = _T_32 & _T_33; // @[HandShaking.scala 218:27]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_18 ? _GEN_22 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_1_valid = _T_18 ? _GEN_23 : out_valid_R_1; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_1_bits_data = _T_18 ? _GEN_16 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_56 = _T_18 & _T_20; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_ready_R_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  out_valid_R_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  value = _RAND_7[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  left_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  left_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  right_R_data = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  right_valid_R = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  state = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  out_data_R = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_4) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_4) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_4) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_4) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_4) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_2) begin
          out_ready_R_1 <= io_Out_1_ready;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_ready_R_1 <= 1'h0;
          end else begin
            if (_T_2) begin
              out_ready_R_1 <= io_Out_1_ready;
            end
          end
        end else begin
          if (_T_2) begin
            out_ready_R_1 <= io_Out_1_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_0 <= _T_25;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      out_valid_R_1 <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          out_valid_R_1 <= _T_26;
        end else begin
          if (_T_2) begin
            out_valid_R_1 <= 1'h0;
          end
        end
      end else begin
        if (_T_2) begin
          out_valid_R_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_7;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_13) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_11;
        end
      end else begin
        left_valid_R <= _GEN_11;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_15) begin
        right_R_data <= 32'h1;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_18) begin
        if (_T_20) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_15;
        end
      end else begin
        right_valid_R <= _GEN_15;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_18) begin
        state <= _GEN_28;
      end else begin
        if (state) begin
          if (_T_34) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_18) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_34) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_56 & _T_28) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] binaryOp_inc105: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ComputeNode_45(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  input         io_Out_0_ready,
  output        io_Out_0_valid,
  output [4:0]  io_Out_0_bits_taskID,
  output [31:0] io_Out_0_bits_data,
  output        io_LeftIO_ready,
  input         io_LeftIO_valid,
  input  [31:0] io_LeftIO_bits_data,
  output        io_RightIO_ready,
  input         io_RightIO_valid
);
  wire [31:0] FU_io_in1; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_in2; // @[ComputeNode.scala 55:18]
  wire [31:0] FU_io_out; // @[ComputeNode.scala 55:18]
  reg [4:0] enable_R_taskID; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_0;
  reg  enable_R_control; // @[HandShaking.scala 167:31]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[HandShaking.scala 168:31]
  reg [31:0] _RAND_2;
  reg  out_ready_R_0; // @[HandShaking.scala 171:46]
  reg [31:0] _RAND_3;
  reg  out_valid_R_0; // @[HandShaking.scala 172:46]
  reg [31:0] _RAND_4;
  wire  _T_1; // @[Decoupled.scala 40:37]
  wire  _T_3; // @[Decoupled.scala 40:37]
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_5;
  wire [14:0] _T_6; // @[Counter.scala 38:22]
  reg [31:0] left_R_data; // @[ComputeNode.scala 47:23]
  reg [31:0] _RAND_6;
  reg  left_valid_R; // @[ComputeNode.scala 48:29]
  reg [31:0] _RAND_7;
  reg [31:0] right_R_data; // @[ComputeNode.scala 51:24]
  reg [31:0] _RAND_8;
  reg  right_valid_R; // @[ComputeNode.scala 52:30]
  reg [31:0] _RAND_9;
  reg  state; // @[ComputeNode.scala 58:22]
  reg [31:0] _RAND_10;
  reg [31:0] out_data_R; // @[ComputeNode.scala 62:27]
  reg [31:0] _RAND_11;
  wire [4:0] taskID; // @[ComputeNode.scala 64:19]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[ComputeNode.scala 74:26]
  wire  _T_14; // @[Decoupled.scala 40:37]
  wire  _GEN_13; // @[ComputeNode.scala 80:27]
  wire  _T_16; // @[Conditional.scala 37:30]
  wire  _T_17; // @[ComputeNode.scala 99:27]
  wire  _T_18; // @[ComputeNode.scala 99:43]
  wire  _T_21; // @[HandShaking.scala 232:72]
  wire  _T_22; // @[ComputeNode.scala 107:17]
  wire  _T_23; // @[ComputeNode.scala 107:17]
  wire [31:0] _T_19_data; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  wire [31:0] _GEN_14; // @[ComputeNode.scala 99:61]
  wire  _GEN_17; // @[ComputeNode.scala 99:61]
  wire  _GEN_21; // @[ComputeNode.scala 99:61]
  wire  _T_26; // @[HandShaking.scala 217:83]
  wire  _GEN_41; // @[ComputeNode.scala 107:17]
  UALU_12 FU ( // @[ComputeNode.scala 55:18]
    .io_in1(FU_io_in1),
    .io_in2(FU_io_in2),
    .io_out(FU_io_out)
  );
  assign _T_1 = io_Out_0_ready & io_Out_0_valid; // @[Decoupled.scala 40:37]
  assign _T_3 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_6 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 64:19]
  assign _T_12 = io_LeftIO_ready & io_LeftIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_12 | left_valid_R; // @[ComputeNode.scala 74:26]
  assign _T_14 = io_RightIO_ready & io_RightIO_valid; // @[Decoupled.scala 40:37]
  assign _GEN_13 = _T_14 | right_valid_R; // @[ComputeNode.scala 80:27]
  assign _T_16 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_17 = enable_valid_R & left_valid_R; // @[ComputeNode.scala 99:27]
  assign _T_18 = _T_17 & right_valid_R; // @[ComputeNode.scala 99:43]
  assign _T_21 = _T_1 ^ 1'h1; // @[HandShaking.scala 232:72]
  assign _T_22 = $unsigned(reset); // @[ComputeNode.scala 107:17]
  assign _T_23 = _T_22 == 1'h0; // @[ComputeNode.scala 107:17]
  assign _T_19_data = FU_io_out; // @[interfaces.scala 305:20 interfaces.scala 306:15]
  assign _GEN_14 = _T_18 ? _T_19_data : out_data_R; // @[ComputeNode.scala 99:61]
  assign _GEN_17 = _T_18 | out_valid_R_0; // @[ComputeNode.scala 99:61]
  assign _GEN_21 = _T_18 | state; // @[ComputeNode.scala 99:61]
  assign _T_26 = out_ready_R_0 | _T_1; // @[HandShaking.scala 217:83]
  assign io_enable_ready = ~ enable_valid_R; // @[HandShaking.scala 191:19]
  assign io_Out_0_valid = _T_16 ? _GEN_17 : out_valid_R_0; // @[HandShaking.scala 180:21 ComputeNode.scala 101:32]
  assign io_Out_0_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_Out_0_bits_data = _T_16 ? _GEN_14 : out_data_R; // @[ComputeNode.scala 92:25 ComputeNode.scala 100:31]
  assign io_LeftIO_ready = ~ left_valid_R; // @[ComputeNode.scala 73:19]
  assign io_RightIO_ready = ~ right_valid_R; // @[ComputeNode.scala 79:20]
  assign FU_io_in1 = left_R_data; // @[ComputeNode.scala 70:13]
  assign FU_io_in2 = right_R_data; // @[ComputeNode.scala 71:13]
  assign _GEN_41 = _T_16 & _T_18; // @[ComputeNode.scala 107:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  enable_R_taskID = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  out_ready_R_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  out_valid_R_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  left_R_data = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  left_valid_R = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  right_R_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  right_valid_R = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  state = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  out_data_R = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_3) begin
        enable_R_taskID <= io_enable_bits_taskID;
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_3) begin
        enable_R_control <= io_enable_bits_control;
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_3) begin
          enable_valid_R <= io_enable_valid;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            enable_valid_R <= 1'h0;
          end else begin
            if (_T_3) begin
              enable_valid_R <= io_enable_valid;
            end
          end
        end else begin
          if (_T_3) begin
            enable_valid_R <= io_enable_valid;
          end
        end
      end
    end
    if (reset) begin
      out_ready_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_1) begin
          out_ready_R_0 <= io_Out_0_ready;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_ready_R_0 <= 1'h0;
          end else begin
            if (_T_1) begin
              out_ready_R_0 <= io_Out_0_ready;
            end
          end
        end else begin
          if (_T_1) begin
            out_ready_R_0 <= io_Out_0_ready;
          end
        end
      end
    end
    if (reset) begin
      out_valid_R_0 <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          out_valid_R_0 <= _T_21;
        end else begin
          if (_T_1) begin
            out_valid_R_0 <= 1'h0;
          end
        end
      end else begin
        if (_T_1) begin
          out_valid_R_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_6;
    end
    if (reset) begin
      left_R_data <= 32'h0;
    end else begin
      if (_T_12) begin
        left_R_data <= io_LeftIO_bits_data;
      end
    end
    if (reset) begin
      left_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          left_valid_R <= 1'h0;
        end else begin
          left_valid_R <= _GEN_9;
        end
      end else begin
        left_valid_R <= _GEN_9;
      end
    end
    if (reset) begin
      right_R_data <= 32'h0;
    end else begin
      if (_T_14) begin
        right_R_data <= 32'h1f;
      end
    end
    if (reset) begin
      right_valid_R <= 1'h0;
    end else begin
      if (_T_16) begin
        if (_T_18) begin
          right_valid_R <= 1'h0;
        end else begin
          right_valid_R <= _GEN_13;
        end
      end else begin
        right_valid_R <= _GEN_13;
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_16) begin
        state <= _GEN_21;
      end else begin
        if (state) begin
          if (_T_26) begin
            state <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      out_data_R <= 32'h0;
    end else begin
      if (_T_16) begin
        if (enable_R_control) begin
          out_data_R <= FU_io_out;
        end else begin
          out_data_R <= 32'h0;
        end
      end else begin
        if (state) begin
          if (_T_26) begin
            out_data_R <= 32'h0;
          end else begin
            if (enable_R_control) begin
              out_data_R <= FU_io_out;
            end else begin
              out_data_R <= 32'h0;
            end
          end
        end else begin
          if (enable_R_control) begin
            out_data_R <= FU_io_out;
          end else begin
            out_data_R <= 32'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_41 & _T_23) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [COMPUTE] icmp_exitcond106: Output fired @ %d, Value: %d (%d + %d)\n",taskID,value,FU_io_out,left_R_data,right_R_data); // @[ComputeNode.scala 107:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CBranchNodeVariable_1(
  input         clock,
  input         reset,
  output        io_enable_ready,
  input         io_enable_valid,
  input  [4:0]  io_enable_bits_taskID,
  input         io_enable_bits_control,
  output        io_CmpIO_ready,
  input         io_CmpIO_valid,
  input  [4:0]  io_CmpIO_bits_taskID,
  input  [31:0] io_CmpIO_bits_data,
  input         io_TrueOutput_0_ready,
  output        io_TrueOutput_0_valid,
  output        io_TrueOutput_0_bits_control,
  input         io_FalseOutput_0_ready,
  output        io_FalseOutput_0_valid,
  output [4:0]  io_FalseOutput_0_bits_taskID,
  output        io_FalseOutput_0_bits_control
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] cmp_R_taskID; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_1;
  reg  cmp_R_control; // @[BranchNode.scala 1193:22]
  reg [31:0] _RAND_2;
  reg  cmp_valid; // @[BranchNode.scala 1194:26]
  reg [31:0] _RAND_3;
  reg [4:0] enable_R_taskID; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_4;
  reg  enable_R_control; // @[BranchNode.scala 1197:25]
  reg [31:0] _RAND_5;
  reg  enable_valid_R; // @[BranchNode.scala 1198:31]
  reg [31:0] _RAND_6;
  reg  output_true_R_control; // @[BranchNode.scala 1204:30]
  reg [31:0] _RAND_7;
  reg  output_true_valid_R_0; // @[BranchNode.scala 1205:54]
  reg [31:0] _RAND_8;
  reg  fire_true_R_0; // @[BranchNode.scala 1206:46]
  reg [31:0] _RAND_9;
  reg [4:0] output_false_R_taskID; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_10;
  reg  output_false_R_control; // @[BranchNode.scala 1208:31]
  reg [31:0] _RAND_11;
  reg  output_false_valid_R_0; // @[BranchNode.scala 1209:56]
  reg [31:0] _RAND_12;
  reg  fire_false_R_0; // @[BranchNode.scala 1210:48]
  reg [31:0] _RAND_13;
  wire [4:0] task_id; // @[BranchNode.scala 1212:33]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_10; // @[BranchNode.scala 1218:44]
  wire  _GEN_3; // @[BranchNode.scala 1217:23]
  wire  _T_12; // @[Decoupled.scala 40:37]
  wire  _GEN_6; // @[BranchNode.scala 1243:24]
  wire  predicate; // @[BranchNode.scala 1249:36]
  wire  true_output; // @[BranchNode.scala 1250:31]
  wire  _T_13; // @[BranchNode.scala 1251:35]
  wire  false_output; // @[BranchNode.scala 1251:32]
  wire  _T_15; // @[Decoupled.scala 40:37]
  wire  _GEN_7; // @[BranchNode.scala 1264:33]
  wire  _GEN_8; // @[BranchNode.scala 1264:33]
  wire  _T_16; // @[Decoupled.scala 40:37]
  wire  _GEN_9; // @[BranchNode.scala 1282:34]
  wire  _GEN_10; // @[BranchNode.scala 1282:34]
  reg  state; // @[BranchNode.scala 1294:22]
  reg [31:0] _RAND_14;
  wire  _T_17; // @[Conditional.scala 37:30]
  wire  _T_18; // @[BranchNode.scala 1300:27]
  wire  _T_20; // @[BranchNode.scala 1310:21]
  wire  _T_21; // @[BranchNode.scala 1310:21]
  wire  _GEN_11; // @[BranchNode.scala 1300:65]
  wire  _GEN_12; // @[BranchNode.scala 1300:65]
  wire  _GEN_13; // @[BranchNode.scala 1300:65]
  wire  _T_27; // @[BranchNode.scala 1334:27]
  wire  _GEN_59; // @[BranchNode.scala 1310:21]
  wire  _GEN_60; // @[BranchNode.scala 1310:21]
  wire  _GEN_62; // @[BranchNode.scala 1324:19]
  wire  _GEN_63; // @[BranchNode.scala 1324:19]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign task_id = enable_R_taskID | cmp_R_taskID; // @[BranchNode.scala 1212:33]
  assign _T_9 = io_CmpIO_ready & io_CmpIO_valid; // @[Decoupled.scala 40:37]
  assign _T_10 = io_CmpIO_bits_data != 32'h0; // @[BranchNode.scala 1218:44]
  assign _GEN_3 = _T_9 | cmp_valid; // @[BranchNode.scala 1217:23]
  assign _T_12 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _GEN_6 = _T_12 | enable_valid_R; // @[BranchNode.scala 1243:24]
  assign predicate = enable_R_control & enable_valid_R; // @[BranchNode.scala 1249:36]
  assign true_output = predicate & cmp_R_control; // @[BranchNode.scala 1250:31]
  assign _T_13 = ~ cmp_R_control; // @[BranchNode.scala 1251:35]
  assign false_output = predicate & _T_13; // @[BranchNode.scala 1251:32]
  assign _T_15 = io_TrueOutput_0_ready & io_TrueOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_7 = _T_15 | fire_true_R_0; // @[BranchNode.scala 1264:33]
  assign _GEN_8 = _T_15 ? 1'h0 : output_true_valid_R_0; // @[BranchNode.scala 1264:33]
  assign _T_16 = io_FalseOutput_0_ready & io_FalseOutput_0_valid; // @[Decoupled.scala 40:37]
  assign _GEN_9 = _T_16 | fire_false_R_0; // @[BranchNode.scala 1282:34]
  assign _GEN_10 = _T_16 ? 1'h0 : output_false_valid_R_0; // @[BranchNode.scala 1282:34]
  assign _T_17 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_18 = enable_valid_R & cmp_valid; // @[BranchNode.scala 1300:27]
  assign _T_20 = $unsigned(reset); // @[BranchNode.scala 1310:21]
  assign _T_21 = _T_20 == 1'h0; // @[BranchNode.scala 1310:21]
  assign _GEN_11 = _T_18 | _GEN_8; // @[BranchNode.scala 1300:65]
  assign _GEN_12 = _T_18 | _GEN_10; // @[BranchNode.scala 1300:65]
  assign _GEN_13 = _T_18 | state; // @[BranchNode.scala 1300:65]
  assign _T_27 = fire_true_R_0 & fire_false_R_0; // @[BranchNode.scala 1334:27]
  assign io_enable_ready = ~ enable_valid_R; // @[BranchNode.scala 1242:19]
  assign io_CmpIO_ready = ~ cmp_valid; // @[BranchNode.scala 1216:18]
  assign io_TrueOutput_0_valid = output_true_valid_R_0; // @[BranchNode.scala 1260:28]
  assign io_TrueOutput_0_bits_control = output_true_R_control; // @[BranchNode.scala 1259:27]
  assign io_FalseOutput_0_valid = output_false_valid_R_0; // @[BranchNode.scala 1278:29]
  assign io_FalseOutput_0_bits_taskID = output_false_R_taskID; // @[BranchNode.scala 1277:28]
  assign io_FalseOutput_0_bits_control = output_false_R_control; // @[BranchNode.scala 1277:28]
  assign _GEN_59 = _T_17 & _T_18; // @[BranchNode.scala 1310:21]
  assign _GEN_60 = _GEN_59 & enable_R_control; // @[BranchNode.scala 1310:21]
  assign _GEN_62 = enable_R_control == 1'h0; // @[BranchNode.scala 1324:19]
  assign _GEN_63 = _GEN_59 & _GEN_62; // @[BranchNode.scala 1324:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cmp_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  cmp_R_control = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  cmp_valid = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  enable_R_taskID = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  enable_R_control = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  enable_valid_R = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  output_true_R_control = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  output_true_valid_R_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  fire_true_R_0 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  output_false_R_taskID = _RAND_10[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  output_false_R_control = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  output_false_valid_R_0 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  fire_false_R_0 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  state = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      cmp_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_taskID <= io_CmpIO_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_taskID <= 5'h0;
          end else begin
            if (_T_9) begin
              cmp_R_taskID <= io_CmpIO_bits_taskID;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_taskID <= io_CmpIO_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      cmp_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_9) begin
          cmp_R_control <= _T_10;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_R_control <= 1'h0;
          end else begin
            if (_T_9) begin
              cmp_R_control <= _T_10;
            end
          end
        end else begin
          if (_T_9) begin
            cmp_R_control <= _T_10;
          end
        end
      end
    end
    if (reset) begin
      cmp_valid <= 1'h0;
    end else begin
      if (_T_17) begin
        cmp_valid <= _GEN_3;
      end else begin
        if (state) begin
          if (_T_27) begin
            cmp_valid <= 1'h0;
          end else begin
            cmp_valid <= _GEN_3;
          end
        end else begin
          cmp_valid <= _GEN_3;
        end
      end
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_taskID <= io_enable_bits_taskID;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_taskID <= 5'h0;
          end else begin
            if (_T_12) begin
              enable_R_taskID <= io_enable_bits_taskID;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end
    end
    if (reset) begin
      enable_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        if (_T_12) begin
          enable_R_control <= io_enable_bits_control;
        end
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_R_control <= 1'h0;
          end else begin
            if (_T_12) begin
              enable_R_control <= io_enable_bits_control;
            end
          end
        end else begin
          if (_T_12) begin
            enable_R_control <= io_enable_bits_control;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_17) begin
        enable_valid_R <= _GEN_6;
      end else begin
        if (state) begin
          if (_T_27) begin
            enable_valid_R <= 1'h0;
          end else begin
            enable_valid_R <= _GEN_6;
          end
        end else begin
          enable_valid_R <= _GEN_6;
        end
      end
    end
    if (reset) begin
      output_true_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_R_control <= true_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_R_control <= 1'h0;
          end else begin
            output_true_R_control <= true_output;
          end
        end else begin
          output_true_R_control <= true_output;
        end
      end
    end
    if (reset) begin
      output_true_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_true_valid_R_0 <= _GEN_11;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_true_valid_R_0 <= 1'h0;
          end else begin
            if (_T_15) begin
              output_true_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_15) begin
            output_true_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_true_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_true_R_0 <= _GEN_7;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_true_R_0 <= 1'h0;
          end else begin
            fire_true_R_0 <= _GEN_7;
          end
        end else begin
          fire_true_R_0 <= _GEN_7;
        end
      end
    end
    if (reset) begin
      output_false_R_taskID <= 5'h0;
    end else begin
      if (_T_17) begin
        output_false_R_taskID <= task_id;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_taskID <= 5'h0;
          end else begin
            output_false_R_taskID <= task_id;
          end
        end else begin
          output_false_R_taskID <= task_id;
        end
      end
    end
    if (reset) begin
      output_false_R_control <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_R_control <= false_output;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_R_control <= 1'h0;
          end else begin
            output_false_R_control <= false_output;
          end
        end else begin
          output_false_R_control <= false_output;
        end
      end
    end
    if (reset) begin
      output_false_valid_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        output_false_valid_R_0 <= _GEN_12;
      end else begin
        if (state) begin
          if (_T_27) begin
            output_false_valid_R_0 <= 1'h0;
          end else begin
            if (_T_16) begin
              output_false_valid_R_0 <= 1'h0;
            end
          end
        end else begin
          if (_T_16) begin
            output_false_valid_R_0 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      fire_false_R_0 <= 1'h0;
    end else begin
      if (_T_17) begin
        fire_false_R_0 <= _GEN_9;
      end else begin
        if (state) begin
          if (_T_27) begin
            fire_false_R_0 <= 1'h0;
          end else begin
            fire_false_R_0 <= _GEN_9;
          end
        end else begin
          fire_false_R_0 <= _GEN_9;
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_17) begin
        state <= _GEN_13;
      end else begin
        if (state) begin
          if (_T_27) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_60 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CBR] br_107: Output fired [T F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1310:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_63 & _T_21) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CBR] br_107: Output fired [F F] @ %d,\n",enable_R_taskID,value); // @[BranchNode.scala 1324:19]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const0: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_1(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const1: Output fired @ %d, Value: %d\n",taskID,value,32'sh2); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_2(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const2: Output fired @ %d, Value: %d\n",taskID,value,32'sh3); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_3(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const3: Output fired @ %d, Value: %d\n",taskID,value,32'sh4); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_4(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const4: Output fired @ %d, Value: %d\n",taskID,value,32'sh5); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_5(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const5: Output fired @ %d, Value: %d\n",taskID,value,32'sh6); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_6(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const6: Output fired @ %d, Value: %d\n",taskID,value,32'sh7); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_7(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const7: Output fired @ %d, Value: %d\n",taskID,value,32'sh8); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_8(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [4:0] io_Out_bits_taskID
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign io_Out_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 126:15]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const8: Output fired @ %d, Value: %d\n",taskID,value,32'sh0); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_9(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const9: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_10(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const10: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_11(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const11: Output fired @ %d, Value: %d\n",taskID,value,32'sh2); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_12(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const12: Output fired @ %d, Value: %d\n",taskID,value,32'sh1f); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_13(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const13: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_14(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const14: Output fired @ %d, Value: %d\n",taskID,value,32'sh1f); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_15(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid,
  output [4:0] io_Out_bits_taskID
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign io_Out_bits_taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 126:15]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const15: Output fired @ %d, Value: %d\n",taskID,value,32'sh0); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_16(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const16: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_17(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const17: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_18(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const18: Output fired @ %d, Value: %d\n",taskID,value,32'sh2); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_19(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const19: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_20(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const20: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_21(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const21: Output fired @ %d, Value: %d\n",taskID,value,32'sh2); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_22(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const22: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_23(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const23: Output fired @ %d, Value: %d\n",taskID,value,32'sh2); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_24(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const24: Output fired @ %d, Value: %d\n",taskID,value,32'sh1); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module ConstFastNode_25(
  input        clock,
  input        reset,
  output       io_enable_ready,
  input        io_enable_valid,
  input  [4:0] io_enable_bits_taskID,
  input        io_Out_ready,
  output       io_Out_valid
);
  reg [14:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire [14:0] _T_2; // @[Counter.scala 38:22]
  reg [4:0] enable_R_taskID; // @[ConstNode.scala 110:25]
  reg [31:0] _RAND_1;
  reg  enable_valid_R; // @[ConstNode.scala 111:31]
  reg [31:0] _RAND_2;
  wire [4:0] taskID; // @[ConstNode.scala 113:19]
  reg  state; // @[ConstNode.scala 132:22]
  reg [31:0] _RAND_3;
  wire  _T_7; // @[Conditional.scala 37:30]
  wire  _T_8; // @[Decoupled.scala 40:37]
  wire  _T_9; // @[Decoupled.scala 40:37]
  wire  _T_11; // @[ConstNode.scala 146:17]
  wire  _T_12; // @[ConstNode.scala 146:17]
  wire  _GEN_5; // @[ConstNode.scala 136:30]
  wire  _GEN_23; // @[ConstNode.scala 146:17]
  assign _T_2 = value + 15'h1; // @[Counter.scala 38:22]
  assign taskID = enable_valid_R ? enable_R_taskID : io_enable_bits_taskID; // @[ConstNode.scala 113:19]
  assign _T_7 = 1'h0 == state; // @[Conditional.scala 37:30]
  assign _T_8 = io_enable_ready & io_enable_valid; // @[Decoupled.scala 40:37]
  assign _T_9 = io_Out_ready & io_Out_valid; // @[Decoupled.scala 40:37]
  assign _T_11 = $unsigned(reset); // @[ConstNode.scala 146:17]
  assign _T_12 = _T_11 == 1'h0; // @[ConstNode.scala 146:17]
  assign _GEN_5 = _T_8 | enable_valid_R; // @[ConstNode.scala 136:30]
  assign io_enable_ready = ~ enable_valid_R; // @[ConstNode.scala 123:19]
  assign io_Out_valid = _T_7 ? _GEN_5 : enable_valid_R; // @[ConstNode.scala 124:16 ConstNode.scala 137:22]
  assign _GEN_23 = _T_7 & _T_8; // @[ConstNode.scala 146:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enable_R_taskID = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enable_valid_R = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end
  always @(posedge clock) begin
    if (reset) begin
      value <= 15'h0;
    end else begin
      value <= _T_2;
    end
    if (reset) begin
      enable_R_taskID <= 5'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_R_taskID <= io_enable_bits_taskID;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_R_taskID <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      enable_valid_R <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (!(_T_9)) begin
            enable_valid_R <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            enable_valid_R <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      state <= 1'h0;
    end else begin
      if (_T_7) begin
        if (_T_8) begin
          if (_T_9) begin
            state <= 1'h0;
          end else begin
            state <= 1'h1;
          end
        end
      end else begin
        if (state) begin
          if (_T_9) begin
            state <= 1'h0;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_23 & _T_12) begin
          $fwrite(32'h80000002,"[LOG] [Extracted_function_conv] [TID->%d] [CONST] const25: Output fired @ %d, Value: %d\n",taskID,value,32'sh1f); // @[ConstNode.scala 146:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module extracted_function_convDF(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [4:0]  io_in_bits_enable_taskID,
  input         io_in_bits_enable_control,
  input         io_in_bits_data_field5_predicate,
  input  [4:0]  io_in_bits_data_field5_taskID,
  input  [31:0] io_in_bits_data_field5_data,
  input         io_in_bits_data_field4_predicate,
  input  [4:0]  io_in_bits_data_field4_taskID,
  input  [31:0] io_in_bits_data_field4_data,
  input         io_in_bits_data_field3_predicate,
  input  [4:0]  io_in_bits_data_field3_taskID,
  input  [31:0] io_in_bits_data_field3_data,
  input         io_in_bits_data_field2_predicate,
  input  [4:0]  io_in_bits_data_field2_taskID,
  input  [31:0] io_in_bits_data_field2_data,
  input         io_in_bits_data_field1_predicate,
  input  [4:0]  io_in_bits_data_field1_taskID,
  input  [31:0] io_in_bits_data_field1_data,
  input         io_in_bits_data_field0_predicate,
  input  [4:0]  io_in_bits_data_field0_taskID,
  input  [31:0] io_in_bits_data_field0_data,
  input         io_MemResp_valid,
  input         io_MemResp_bits_valid,
  input  [31:0] io_MemResp_bits_data,
  input  [7:0]  io_MemResp_bits_tag,
  input         io_MemResp_bits_iswrite,
  input  [31:0] io_MemResp_bits_tile,
  input         io_MemReq_ready,
  output        io_MemReq_valid,
  output [31:0] io_MemReq_bits_addr,
  output [31:0] io_MemReq_bits_data,
  output [3:0]  io_MemReq_bits_mask,
  output [7:0]  io_MemReq_bits_tag,
  output [4:0]  io_MemReq_bits_taskID,
  output        io_MemReq_bits_iswrite,
  output [31:0] io_MemReq_bits_tile,
  input         io_out_ready,
  output        io_out_valid,
  output [4:0]  io_out_bits_enable_taskID,
  output        io_out_bits_enable_control
);
  wire  MemCtrl_clock; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_reset; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_0_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_0_valid; // @[extracted_function_conv.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_0_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_0_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_0_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_1_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_1_valid; // @[extracted_function_conv.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_1_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_1_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_1_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_2_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_2_valid; // @[extracted_function_conv.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_2_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_2_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_2_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_3_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_3_valid; // @[extracted_function_conv.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_3_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_3_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_3_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_4_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_4_valid; // @[extracted_function_conv.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_4_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_4_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_4_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_5_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_5_valid; // @[extracted_function_conv.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_5_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_5_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_5_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_6_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_6_valid; // @[extracted_function_conv.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_6_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_6_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_6_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_7_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_7_valid; // @[extracted_function_conv.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_7_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_7_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_7_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_8_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteIn_8_valid; // @[extracted_function_conv.scala 45:23]
  wire [21:0] MemCtrl_io_WriteIn_8_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_WriteIn_8_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_WriteIn_8_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteOut_0_valid; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteOut_1_valid; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteOut_2_valid; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteOut_3_valid; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteOut_4_valid; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteOut_5_valid; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteOut_6_valid; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteOut_7_valid; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_WriteOut_8_valid; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_0_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_0_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_0_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_0_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_1_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_1_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_1_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_1_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_2_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_2_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_2_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_2_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_3_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_3_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_3_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_3_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_4_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_4_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_4_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_4_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_5_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_5_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_5_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_5_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_6_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_6_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_6_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_6_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_7_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_7_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_7_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_7_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_8_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_8_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_8_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_8_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_9_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_9_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_9_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_9_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_10_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_10_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_10_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_10_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_11_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_11_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_11_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_11_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_12_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_12_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_12_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_12_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_13_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_13_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_13_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_13_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_14_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_14_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_14_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_14_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_15_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_15_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_15_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_15_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_16_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_16_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_16_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_16_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_17_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_17_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_17_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_17_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_18_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadIn_18_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadIn_18_bits_address; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_ReadIn_18_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_0_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_0_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_1_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_1_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_2_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_2_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_3_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_3_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_4_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_4_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_5_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_5_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_6_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_6_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_7_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_7_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_8_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_8_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_9_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_9_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_10_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_10_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_11_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_11_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_12_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_12_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_13_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_13_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_14_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_14_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_15_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_15_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_16_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_16_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_17_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_17_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_ReadOut_18_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_ReadOut_18_data; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_MemResp_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_MemResp_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [7:0] MemCtrl_io_MemResp_bits_tag; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_MemResp_bits_iswrite; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_MemReq_ready; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_MemReq_valid; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_MemReq_bits_addr; // @[extracted_function_conv.scala 45:23]
  wire [31:0] MemCtrl_io_MemReq_bits_data; // @[extracted_function_conv.scala 45:23]
  wire [3:0] MemCtrl_io_MemReq_bits_mask; // @[extracted_function_conv.scala 45:23]
  wire [7:0] MemCtrl_io_MemReq_bits_tag; // @[extracted_function_conv.scala 45:23]
  wire [4:0] MemCtrl_io_MemReq_bits_taskID; // @[extracted_function_conv.scala 45:23]
  wire  MemCtrl_io_MemReq_bits_iswrite; // @[extracted_function_conv.scala 45:23]
  wire  InputSplitter_clock; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_reset; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_In_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_In_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_enable_taskID; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_In_bits_enable_control; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field5_data; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field4_data; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field3_data; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_data_field2_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field2_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_In_bits_data_field1_predicate; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_data_field1_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field1_data; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_In_bits_data_field0_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_In_bits_data_field0_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_enable_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_enable_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_enable_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_enable_bits_control; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field5_0_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field5_0_valid; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field5_0_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field5_1_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field5_1_valid; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field5_1_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field4_0_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field4_0_valid; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field4_0_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field3_0_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field3_0_valid; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field3_0_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field2_0_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field2_0_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field2_0_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field2_0_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_0_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_0_valid; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_0_bits_predicate; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_0_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_0_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_1_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_1_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_1_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_1_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_2_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_2_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_2_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_2_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_3_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_3_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_3_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_3_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_4_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_4_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_4_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_4_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_5_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_5_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_5_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_5_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_6_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_6_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_6_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_6_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_7_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_7_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_7_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_7_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_8_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field1_8_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field1_8_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field1_8_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field0_0_ready; // @[extracted_function_conv.scala 53:29]
  wire  InputSplitter_io_Out_data_field0_0_valid; // @[extracted_function_conv.scala 53:29]
  wire [4:0] InputSplitter_io_Out_data_field0_0_bits_taskID; // @[extracted_function_conv.scala 53:29]
  wire [31:0] InputSplitter_io_Out_data_field0_0_bits_data; // @[extracted_function_conv.scala 53:29]
  wire  Loop_0_clock; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_reset; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_enable_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_enable_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_enable_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_enable_bits_control; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_1_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_1_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_1_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_2_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_2_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_2_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_3_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_3_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_3_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_4_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_4_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_4_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_4_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_4_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_5_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_5_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_5_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_6_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_6_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_6_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_6_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_6_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_7_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_7_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_7_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_7_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_7_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_8_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_8_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_8_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_8_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_8_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_9_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_9_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_9_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_9_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_9_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_10_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_10_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_10_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_10_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_11_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_11_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_11_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_11_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_12_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_12_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_12_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_12_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_12_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_13_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_13_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_13_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_13_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_13_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_14_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_14_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_14_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_14_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_14_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_15_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_15_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_InLiveIn_15_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_InLiveIn_15_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_InLiveIn_15_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field15_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field15_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field15_0_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field15_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field15_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field14_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field14_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field14_0_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field14_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field14_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field13_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field13_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field13_0_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field13_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field13_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field12_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field12_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field12_0_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field12_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field12_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field11_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field11_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field11_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field11_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field10_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field10_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_1_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_1_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field10_1_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field10_1_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_2_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_2_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field10_2_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field10_2_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_3_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_3_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field10_3_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field10_3_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_4_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_4_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field10_4_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field10_4_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_5_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_5_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field10_5_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field10_5_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_6_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_6_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field10_6_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field10_6_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_7_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_7_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field10_7_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field10_7_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_8_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field10_8_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field10_8_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field10_8_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field9_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field9_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field9_0_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field9_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field9_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field8_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field8_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field8_0_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field7_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field7_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field7_0_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field7_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field6_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field6_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field6_0_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field6_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field5_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field5_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field4_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field4_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field4_0_bits_predicate; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field3_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field3_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field2_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field2_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field1_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field1_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field0_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_OutLiveIn_field0_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_activate_loop_start_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_activate_loop_start_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_activate_loop_start_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_activate_loop_start_bits_control; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_activate_loop_back_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_activate_loop_back_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_activate_loop_back_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_activate_loop_back_bits_control; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_loopBack_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_loopBack_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_loopBack_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_loopBack_0_bits_control; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_loopFinish_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_loopFinish_0_valid; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_loopFinish_0_bits_control; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_CarryDepenIn_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_CarryDepenIn_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_CarryDepenIn_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_CarryDepenIn_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_CarryDepenOut_field0_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_CarryDepenOut_field0_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire [31:0] Loop_0_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_loopExit_0_ready; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_loopExit_0_valid; // @[extracted_function_conv.scala 62:22]
  wire [4:0] Loop_0_io_loopExit_0_bits_taskID; // @[extracted_function_conv.scala 62:22]
  wire  Loop_0_io_loopExit_0_bits_control; // @[extracted_function_conv.scala 62:22]
  wire  Loop_1_clock; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_reset; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_enable_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_enable_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_enable_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_enable_bits_control; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_0_valid; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_1_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_1_valid; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_1_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_2_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_2_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_2_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_2_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_3_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_3_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_3_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_3_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_3_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_4_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_4_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_4_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_4_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_5_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_5_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_5_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_5_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_5_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_6_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_6_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_6_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_6_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_6_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_7_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_7_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_7_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_7_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_7_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_8_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_8_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_8_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_8_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_8_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_9_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_9_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_9_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_9_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_9_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_10_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_10_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_10_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_10_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_10_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_11_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_11_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_11_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_11_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_11_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_12_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_12_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_InLiveIn_12_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_InLiveIn_12_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_InLiveIn_12_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field12_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field12_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field12_0_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field12_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field12_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field11_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field11_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field11_0_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field11_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field11_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field10_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field10_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field10_0_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field10_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field10_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field9_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field9_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field9_0_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field9_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field9_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field8_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field8_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field8_0_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field7_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field7_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field7_0_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field7_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field6_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field6_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field6_0_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field6_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field5_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field5_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field5_0_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field5_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field4_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field4_0_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field3_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field3_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field3_0_bits_predicate; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field3_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field2_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field2_0_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_OutLiveIn_field2_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_0_valid; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_1_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_1_valid; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field1_1_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_2_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field1_2_valid; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field1_2_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_0_valid; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_1_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_1_valid; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field0_1_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_2_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_OutLiveIn_field0_2_valid; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_OutLiveIn_field0_2_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_activate_loop_start_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_activate_loop_start_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_activate_loop_start_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_activate_loop_start_bits_control; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_activate_loop_back_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_activate_loop_back_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_activate_loop_back_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_activate_loop_back_bits_control; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_loopBack_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_loopBack_0_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_loopBack_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_loopBack_0_bits_control; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_loopFinish_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_loopFinish_0_valid; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_loopFinish_0_bits_control; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_CarryDepenIn_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_CarryDepenIn_0_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_CarryDepenIn_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_CarryDepenIn_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_CarryDepenOut_field0_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_CarryDepenOut_field0_0_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire [31:0] Loop_1_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_loopExit_0_ready; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_loopExit_0_valid; // @[extracted_function_conv.scala 64:22]
  wire [4:0] Loop_1_io_loopExit_0_bits_taskID; // @[extracted_function_conv.scala 64:22]
  wire  Loop_1_io_loopExit_0_bits_control; // @[extracted_function_conv.scala 64:22]
  wire  bb_entry0_clock; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_reset; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_predicateIn_0_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_predicateIn_0_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_predicateIn_0_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_predicateIn_0_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_0_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_0_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_1_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_1_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_2_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_2_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_3_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_3_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_4_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_4_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_5_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_5_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_5_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_6_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_6_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_6_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_7_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_7_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_7_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_8_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_8_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_8_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_8_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_9_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_9_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_9_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_9_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_10_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_10_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_10_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_10_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_11_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_11_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_11_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_11_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_12_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_12_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_12_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_12_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_13_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_13_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_13_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_13_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_14_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_14_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_14_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_14_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_15_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_15_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_15_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_15_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_16_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_16_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_16_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_16_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_17_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_17_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_17_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_17_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_18_ready; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_18_valid; // @[extracted_function_conv.scala 72:25]
  wire [4:0] bb_entry0_io_Out_18_bits_taskID; // @[extracted_function_conv.scala 72:25]
  wire  bb_entry0_io_Out_18_bits_control; // @[extracted_function_conv.scala 72:25]
  wire  bb_for_cond_cleanup1_clock; // @[extracted_function_conv.scala 74:36]
  wire  bb_for_cond_cleanup1_reset; // @[extracted_function_conv.scala 74:36]
  wire  bb_for_cond_cleanup1_io_predicateIn_0_ready; // @[extracted_function_conv.scala 74:36]
  wire  bb_for_cond_cleanup1_io_predicateIn_0_valid; // @[extracted_function_conv.scala 74:36]
  wire [4:0] bb_for_cond_cleanup1_io_predicateIn_0_bits_taskID; // @[extracted_function_conv.scala 74:36]
  wire  bb_for_cond_cleanup1_io_predicateIn_0_bits_control; // @[extracted_function_conv.scala 74:36]
  wire  bb_for_cond_cleanup1_io_Out_0_ready; // @[extracted_function_conv.scala 74:36]
  wire  bb_for_cond_cleanup1_io_Out_0_valid; // @[extracted_function_conv.scala 74:36]
  wire [4:0] bb_for_cond_cleanup1_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 74:36]
  wire  bb_for_cond_cleanup1_io_Out_0_bits_control; // @[extracted_function_conv.scala 74:36]
  wire  bb_for_body2_clock; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_reset; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_MaskBB_0_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_MaskBB_0_valid; // @[extracted_function_conv.scala 76:28]
  wire [1:0] bb_for_body2_io_MaskBB_0_bits; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_0_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_0_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_1_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_1_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_2_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_2_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_3_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_3_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_4_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_4_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_5_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_5_valid; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_5_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_6_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_6_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_6_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_6_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_7_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_7_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_7_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_7_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_8_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_8_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_8_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_8_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_9_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_9_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_9_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_9_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_10_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_10_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_10_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_10_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_11_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_11_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_11_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_11_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_12_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_12_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_12_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_12_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_13_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_13_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_13_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_13_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_14_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_14_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_14_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_14_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_15_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_15_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_Out_15_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_Out_15_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_predicateIn_0_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_predicateIn_0_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_predicateIn_0_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_predicateIn_0_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_predicateIn_1_ready; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_predicateIn_1_valid; // @[extracted_function_conv.scala 76:28]
  wire [4:0] bb_for_body2_io_predicateIn_1_bits_taskID; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_body2_io_predicateIn_1_bits_control; // @[extracted_function_conv.scala 76:28]
  wire  bb_for_cond_cleanup113_clock; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_reset; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_predicateIn_0_ready; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_predicateIn_0_valid; // @[extracted_function_conv.scala 78:38]
  wire [4:0] bb_for_cond_cleanup113_io_predicateIn_0_bits_taskID; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_predicateIn_0_bits_control; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_0_ready; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_0_valid; // @[extracted_function_conv.scala 78:38]
  wire [4:0] bb_for_cond_cleanup113_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_1_ready; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_1_valid; // @[extracted_function_conv.scala 78:38]
  wire [4:0] bb_for_cond_cleanup113_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_2_ready; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_2_valid; // @[extracted_function_conv.scala 78:38]
  wire [4:0] bb_for_cond_cleanup113_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_2_bits_control; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_3_ready; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_3_valid; // @[extracted_function_conv.scala 78:38]
  wire [4:0] bb_for_cond_cleanup113_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_3_bits_control; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_4_ready; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_4_valid; // @[extracted_function_conv.scala 78:38]
  wire [4:0] bb_for_cond_cleanup113_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_cond_cleanup113_io_Out_4_bits_control; // @[extracted_function_conv.scala 78:38]
  wire  bb_for_body124_clock; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_reset; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_MaskBB_0_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_MaskBB_0_valid; // @[extracted_function_conv.scala 80:30]
  wire [1:0] bb_for_body124_io_MaskBB_0_bits; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_0_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_0_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_1_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_1_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_2_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_2_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_3_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_3_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_4_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_4_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_5_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_5_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_5_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_6_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_6_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_6_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_7_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_7_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_7_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_8_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_8_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_8_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_9_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_9_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_9_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_10_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_10_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_10_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_11_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_11_valid; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_11_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_12_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_12_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_12_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_12_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_13_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_13_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_13_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_13_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_14_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_14_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_14_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_14_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_15_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_15_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_15_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_15_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_16_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_16_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_16_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_16_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_17_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_17_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_17_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_17_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_18_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_18_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_18_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_18_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_19_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_19_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_19_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_19_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_20_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_20_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_20_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_20_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_21_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_21_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_21_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_22_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_22_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_22_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_22_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_23_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_23_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_23_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_23_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_24_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_24_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_24_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_24_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_25_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_25_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_25_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_25_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_26_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_26_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_26_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_26_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_27_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_27_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_27_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_27_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_28_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_28_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_28_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_28_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_29_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_29_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_29_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_30_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_30_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_30_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_30_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_31_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_31_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_31_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_31_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_32_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_32_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_32_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_32_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_33_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_33_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_33_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_33_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_34_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_34_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_34_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_34_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_35_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_35_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_35_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_35_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_36_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_36_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_36_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_36_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_37_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_37_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_37_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_38_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_38_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_38_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_38_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_39_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_39_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_39_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_39_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_40_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_40_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_40_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_40_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_41_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_41_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_41_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_41_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_42_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_42_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_42_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_42_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_43_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_43_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_43_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_43_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_44_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_44_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_44_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_44_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_45_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_45_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_45_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_45_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_46_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_46_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_46_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_47_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_47_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_47_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_47_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_48_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_48_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_48_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_48_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_49_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_49_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_49_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_49_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_50_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_50_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_50_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_50_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_51_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_51_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_51_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_51_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_52_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_52_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_52_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_52_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_53_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_53_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_53_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_53_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_54_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_54_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_54_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_55_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_55_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_55_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_55_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_56_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_56_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_56_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_56_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_57_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_57_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_57_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_57_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_58_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_58_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_58_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_58_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_59_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_59_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_59_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_59_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_60_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_60_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_60_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_60_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_61_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_61_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_61_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_61_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_62_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_62_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_62_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_63_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_63_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_63_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_63_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_64_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_64_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_64_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_64_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_65_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_65_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_65_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_65_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_66_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_66_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_66_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_66_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_67_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_67_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_67_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_67_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_68_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_68_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_68_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_68_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_69_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_69_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_69_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_69_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_70_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_70_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_70_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_71_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_71_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_71_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_71_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_72_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_72_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_72_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_72_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_73_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_73_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_73_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_73_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_74_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_74_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_74_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_74_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_75_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_75_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_75_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_75_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_76_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_76_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_76_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_76_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_77_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_77_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_77_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_77_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_78_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_78_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_78_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_79_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_79_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_79_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_79_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_80_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_80_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_80_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_80_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_81_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_81_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_81_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_81_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_82_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_82_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_82_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_82_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_83_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_83_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_83_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_83_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_84_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_84_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_84_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_84_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_85_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_85_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_85_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_85_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_86_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_86_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_86_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_87_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_87_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_87_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_87_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_88_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_88_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_88_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_88_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_89_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_89_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_89_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_89_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_90_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_90_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_90_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_90_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_91_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_91_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_91_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_91_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_92_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_92_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_Out_92_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_Out_92_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_predicateIn_0_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_predicateIn_0_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_predicateIn_0_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_predicateIn_0_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_predicateIn_1_ready; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_predicateIn_1_valid; // @[extracted_function_conv.scala 80:30]
  wire [4:0] bb_for_body124_io_predicateIn_1_bits_taskID; // @[extracted_function_conv.scala 80:30]
  wire  bb_for_body124_io_predicateIn_1_bits_control; // @[extracted_function_conv.scala 80:30]
  wire  binaryOp_mul0_clock; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_reset; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_io_enable_ready; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_io_enable_valid; // @[extracted_function_conv.scala 89:29]
  wire [4:0] binaryOp_mul0_io_enable_bits_taskID; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_io_enable_bits_control; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_io_Out_0_ready; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_io_Out_0_valid; // @[extracted_function_conv.scala 89:29]
  wire [31:0] binaryOp_mul0_io_Out_0_bits_data; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_io_LeftIO_ready; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_io_LeftIO_valid; // @[extracted_function_conv.scala 89:29]
  wire [31:0] binaryOp_mul0_io_LeftIO_bits_data; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_io_RightIO_ready; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_mul0_io_RightIO_valid; // @[extracted_function_conv.scala 89:29]
  wire [31:0] binaryOp_mul0_io_RightIO_bits_data; // @[extracted_function_conv.scala 89:29]
  wire  binaryOp_add1_clock; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_reset; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_io_enable_ready; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_io_enable_valid; // @[extracted_function_conv.scala 92:29]
  wire [4:0] binaryOp_add1_io_enable_bits_taskID; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_io_enable_bits_control; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_io_Out_0_ready; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_io_Out_0_valid; // @[extracted_function_conv.scala 92:29]
  wire [31:0] binaryOp_add1_io_Out_0_bits_data; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_io_LeftIO_ready; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_io_LeftIO_valid; // @[extracted_function_conv.scala 92:29]
  wire [31:0] binaryOp_add1_io_LeftIO_bits_data; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_io_RightIO_ready; // @[extracted_function_conv.scala 92:29]
  wire  binaryOp_add1_io_RightIO_valid; // @[extracted_function_conv.scala 92:29]
  wire [31:0] binaryOp_add1_io_RightIO_bits_data; // @[extracted_function_conv.scala 92:29]
  wire  Gep_arrayidx252_clock; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_reset; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_enable_ready; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_enable_valid; // @[extracted_function_conv.scala 95:31]
  wire [4:0] Gep_arrayidx252_io_enable_bits_taskID; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_enable_bits_control; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_Out_0_ready; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_Out_0_valid; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 95:31]
  wire [4:0] Gep_arrayidx252_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 95:31]
  wire [31:0] Gep_arrayidx252_io_Out_0_bits_data; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_baseAddress_ready; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_baseAddress_valid; // @[extracted_function_conv.scala 95:31]
  wire [4:0] Gep_arrayidx252_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 95:31]
  wire [31:0] Gep_arrayidx252_io_baseAddress_bits_data; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_idx_0_ready; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx252_io_idx_0_valid; // @[extracted_function_conv.scala 95:31]
  wire  Gep_arrayidx383_clock; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_reset; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_enable_ready; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_enable_valid; // @[extracted_function_conv.scala 98:31]
  wire [4:0] Gep_arrayidx383_io_enable_bits_taskID; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_enable_bits_control; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_Out_0_ready; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_Out_0_valid; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 98:31]
  wire [4:0] Gep_arrayidx383_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 98:31]
  wire [31:0] Gep_arrayidx383_io_Out_0_bits_data; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_baseAddress_ready; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_baseAddress_valid; // @[extracted_function_conv.scala 98:31]
  wire [4:0] Gep_arrayidx383_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 98:31]
  wire [31:0] Gep_arrayidx383_io_baseAddress_bits_data; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_idx_0_ready; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx383_io_idx_0_valid; // @[extracted_function_conv.scala 98:31]
  wire  Gep_arrayidx514_clock; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_reset; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_enable_ready; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_enable_valid; // @[extracted_function_conv.scala 101:31]
  wire [4:0] Gep_arrayidx514_io_enable_bits_taskID; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_enable_bits_control; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_Out_0_ready; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_Out_0_valid; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 101:31]
  wire [4:0] Gep_arrayidx514_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 101:31]
  wire [31:0] Gep_arrayidx514_io_Out_0_bits_data; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_baseAddress_ready; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_baseAddress_valid; // @[extracted_function_conv.scala 101:31]
  wire [4:0] Gep_arrayidx514_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 101:31]
  wire [31:0] Gep_arrayidx514_io_baseAddress_bits_data; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_idx_0_ready; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx514_io_idx_0_valid; // @[extracted_function_conv.scala 101:31]
  wire  Gep_arrayidx625_clock; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_reset; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_enable_ready; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_enable_valid; // @[extracted_function_conv.scala 104:31]
  wire [4:0] Gep_arrayidx625_io_enable_bits_taskID; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_enable_bits_control; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_Out_0_ready; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_Out_0_valid; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 104:31]
  wire [4:0] Gep_arrayidx625_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 104:31]
  wire [31:0] Gep_arrayidx625_io_Out_0_bits_data; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_baseAddress_ready; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_baseAddress_valid; // @[extracted_function_conv.scala 104:31]
  wire [4:0] Gep_arrayidx625_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 104:31]
  wire [31:0] Gep_arrayidx625_io_baseAddress_bits_data; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_idx_0_ready; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx625_io_idx_0_valid; // @[extracted_function_conv.scala 104:31]
  wire  Gep_arrayidx746_clock; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_reset; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_enable_ready; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_enable_valid; // @[extracted_function_conv.scala 107:31]
  wire [4:0] Gep_arrayidx746_io_enable_bits_taskID; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_enable_bits_control; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_Out_0_ready; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_Out_0_valid; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 107:31]
  wire [4:0] Gep_arrayidx746_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 107:31]
  wire [31:0] Gep_arrayidx746_io_Out_0_bits_data; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_baseAddress_ready; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_baseAddress_valid; // @[extracted_function_conv.scala 107:31]
  wire [4:0] Gep_arrayidx746_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 107:31]
  wire [31:0] Gep_arrayidx746_io_baseAddress_bits_data; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_idx_0_ready; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx746_io_idx_0_valid; // @[extracted_function_conv.scala 107:31]
  wire  Gep_arrayidx867_clock; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_reset; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_enable_ready; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_enable_valid; // @[extracted_function_conv.scala 110:31]
  wire [4:0] Gep_arrayidx867_io_enable_bits_taskID; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_enable_bits_control; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_Out_0_ready; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_Out_0_valid; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 110:31]
  wire [4:0] Gep_arrayidx867_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 110:31]
  wire [31:0] Gep_arrayidx867_io_Out_0_bits_data; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_baseAddress_ready; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_baseAddress_valid; // @[extracted_function_conv.scala 110:31]
  wire [4:0] Gep_arrayidx867_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 110:31]
  wire [31:0] Gep_arrayidx867_io_baseAddress_bits_data; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_idx_0_ready; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx867_io_idx_0_valid; // @[extracted_function_conv.scala 110:31]
  wire  Gep_arrayidx978_clock; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_reset; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_enable_ready; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_enable_valid; // @[extracted_function_conv.scala 113:31]
  wire [4:0] Gep_arrayidx978_io_enable_bits_taskID; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_enable_bits_control; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_Out_0_ready; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_Out_0_valid; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 113:31]
  wire [4:0] Gep_arrayidx978_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 113:31]
  wire [31:0] Gep_arrayidx978_io_Out_0_bits_data; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_baseAddress_ready; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_baseAddress_valid; // @[extracted_function_conv.scala 113:31]
  wire [4:0] Gep_arrayidx978_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 113:31]
  wire [31:0] Gep_arrayidx978_io_baseAddress_bits_data; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_idx_0_ready; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx978_io_idx_0_valid; // @[extracted_function_conv.scala 113:31]
  wire  Gep_arrayidx1099_clock; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_reset; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_enable_ready; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_enable_valid; // @[extracted_function_conv.scala 116:32]
  wire [4:0] Gep_arrayidx1099_io_enable_bits_taskID; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_enable_bits_control; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_Out_0_ready; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_Out_0_valid; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 116:32]
  wire [4:0] Gep_arrayidx1099_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 116:32]
  wire [31:0] Gep_arrayidx1099_io_Out_0_bits_data; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_baseAddress_ready; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_baseAddress_valid; // @[extracted_function_conv.scala 116:32]
  wire [4:0] Gep_arrayidx1099_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 116:32]
  wire [31:0] Gep_arrayidx1099_io_baseAddress_bits_data; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_idx_0_ready; // @[extracted_function_conv.scala 116:32]
  wire  Gep_arrayidx1099_io_idx_0_valid; // @[extracted_function_conv.scala 116:32]
  wire  br_10_clock; // @[extracted_function_conv.scala 119:21]
  wire  br_10_reset; // @[extracted_function_conv.scala 119:21]
  wire  br_10_io_enable_ready; // @[extracted_function_conv.scala 119:21]
  wire  br_10_io_enable_valid; // @[extracted_function_conv.scala 119:21]
  wire [4:0] br_10_io_enable_bits_taskID; // @[extracted_function_conv.scala 119:21]
  wire  br_10_io_enable_bits_control; // @[extracted_function_conv.scala 119:21]
  wire  br_10_io_Out_0_ready; // @[extracted_function_conv.scala 119:21]
  wire  br_10_io_Out_0_valid; // @[extracted_function_conv.scala 119:21]
  wire [4:0] br_10_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 119:21]
  wire  br_10_io_Out_0_bits_control; // @[extracted_function_conv.scala 119:21]
  wire  ret_11_clock; // @[extracted_function_conv.scala 122:22]
  wire  ret_11_reset; // @[extracted_function_conv.scala 122:22]
  wire  ret_11_io_In_enable_ready; // @[extracted_function_conv.scala 122:22]
  wire  ret_11_io_In_enable_valid; // @[extracted_function_conv.scala 122:22]
  wire [4:0] ret_11_io_In_enable_bits_taskID; // @[extracted_function_conv.scala 122:22]
  wire  ret_11_io_In_enable_bits_control; // @[extracted_function_conv.scala 122:22]
  wire  ret_11_io_Out_ready; // @[extracted_function_conv.scala 122:22]
  wire  ret_11_io_Out_valid; // @[extracted_function_conv.scala 122:22]
  wire [4:0] ret_11_io_Out_bits_enable_taskID; // @[extracted_function_conv.scala 122:22]
  wire  ret_11_io_Out_bits_enable_control; // @[extracted_function_conv.scala 122:22]
  wire  phi_conv_s1_y_031312_clock; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_reset; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_enable_ready; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_enable_valid; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_enable_bits_control; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_InData_0_ready; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_InData_0_valid; // @[extracted_function_conv.scala 125:36]
  wire [4:0] phi_conv_s1_y_031312_io_InData_0_bits_taskID; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_InData_1_ready; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_InData_1_valid; // @[extracted_function_conv.scala 125:36]
  wire [4:0] phi_conv_s1_y_031312_io_InData_1_bits_taskID; // @[extracted_function_conv.scala 125:36]
  wire [31:0] phi_conv_s1_y_031312_io_InData_1_bits_data; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Mask_ready; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Mask_valid; // @[extracted_function_conv.scala 125:36]
  wire [1:0] phi_conv_s1_y_031312_io_Mask_bits; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Out_0_ready; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Out_0_valid; // @[extracted_function_conv.scala 125:36]
  wire [31:0] phi_conv_s1_y_031312_io_Out_0_bits_data; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Out_1_ready; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Out_1_valid; // @[extracted_function_conv.scala 125:36]
  wire [31:0] phi_conv_s1_y_031312_io_Out_1_bits_data; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Out_2_ready; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Out_2_valid; // @[extracted_function_conv.scala 125:36]
  wire [31:0] phi_conv_s1_y_031312_io_Out_2_bits_data; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Out_3_ready; // @[extracted_function_conv.scala 125:36]
  wire  phi_conv_s1_y_031312_io_Out_3_valid; // @[extracted_function_conv.scala 125:36]
  wire [31:0] phi_conv_s1_y_031312_io_Out_3_bits_data; // @[extracted_function_conv.scala 125:36]
  wire  binaryOp_mul113_clock; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_reset; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_enable_ready; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_enable_valid; // @[extracted_function_conv.scala 128:31]
  wire [4:0] binaryOp_mul113_io_enable_bits_taskID; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_enable_bits_control; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_Out_0_ready; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_Out_0_valid; // @[extracted_function_conv.scala 128:31]
  wire [31:0] binaryOp_mul113_io_Out_0_bits_data; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_Out_1_ready; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_Out_1_valid; // @[extracted_function_conv.scala 128:31]
  wire [31:0] binaryOp_mul113_io_Out_1_bits_data; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_LeftIO_ready; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_LeftIO_valid; // @[extracted_function_conv.scala 128:31]
  wire [31:0] binaryOp_mul113_io_LeftIO_bits_data; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_RightIO_ready; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_mul113_io_RightIO_valid; // @[extracted_function_conv.scala 128:31]
  wire  binaryOp_add214_clock; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_reset; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_io_enable_ready; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_io_enable_valid; // @[extracted_function_conv.scala 131:31]
  wire [4:0] binaryOp_add214_io_enable_bits_taskID; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_io_enable_bits_control; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_io_Out_0_ready; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_io_Out_0_valid; // @[extracted_function_conv.scala 131:31]
  wire [31:0] binaryOp_add214_io_Out_0_bits_data; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_io_LeftIO_ready; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_io_LeftIO_valid; // @[extracted_function_conv.scala 131:31]
  wire [31:0] binaryOp_add214_io_LeftIO_bits_data; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_io_RightIO_ready; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_add214_io_RightIO_valid; // @[extracted_function_conv.scala 131:31]
  wire  binaryOp_mul315_clock; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_reset; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_io_enable_ready; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_io_enable_valid; // @[extracted_function_conv.scala 134:31]
  wire [4:0] binaryOp_mul315_io_enable_bits_taskID; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_io_enable_bits_control; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_io_Out_0_ready; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_io_Out_0_valid; // @[extracted_function_conv.scala 134:31]
  wire [31:0] binaryOp_mul315_io_Out_0_bits_data; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_io_LeftIO_ready; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_io_LeftIO_valid; // @[extracted_function_conv.scala 134:31]
  wire [31:0] binaryOp_mul315_io_LeftIO_bits_data; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_io_RightIO_ready; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_mul315_io_RightIO_valid; // @[extracted_function_conv.scala 134:31]
  wire [31:0] binaryOp_mul315_io_RightIO_bits_data; // @[extracted_function_conv.scala 134:31]
  wire  binaryOp_sub16_clock; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_reset; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_io_enable_ready; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_io_enable_valid; // @[extracted_function_conv.scala 137:30]
  wire [4:0] binaryOp_sub16_io_enable_bits_taskID; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_io_enable_bits_control; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_io_Out_0_ready; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_io_Out_0_valid; // @[extracted_function_conv.scala 137:30]
  wire [31:0] binaryOp_sub16_io_Out_0_bits_data; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_io_LeftIO_ready; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_io_LeftIO_valid; // @[extracted_function_conv.scala 137:30]
  wire [31:0] binaryOp_sub16_io_LeftIO_bits_data; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_io_RightIO_ready; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_sub16_io_RightIO_valid; // @[extracted_function_conv.scala 137:30]
  wire [31:0] binaryOp_sub16_io_RightIO_bits_data; // @[extracted_function_conv.scala 137:30]
  wire  binaryOp_add417_clock; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_reset; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_io_enable_ready; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_io_enable_valid; // @[extracted_function_conv.scala 140:31]
  wire [4:0] binaryOp_add417_io_enable_bits_taskID; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_io_enable_bits_control; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_io_Out_0_ready; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_io_Out_0_valid; // @[extracted_function_conv.scala 140:31]
  wire [31:0] binaryOp_add417_io_Out_0_bits_data; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_io_LeftIO_ready; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_io_LeftIO_valid; // @[extracted_function_conv.scala 140:31]
  wire [31:0] binaryOp_add417_io_LeftIO_bits_data; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_io_RightIO_ready; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_add417_io_RightIO_valid; // @[extracted_function_conv.scala 140:31]
  wire  binaryOp_mul518_clock; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_reset; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_io_enable_ready; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_io_enable_valid; // @[extracted_function_conv.scala 143:31]
  wire [4:0] binaryOp_mul518_io_enable_bits_taskID; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_io_enable_bits_control; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_io_Out_0_ready; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_io_Out_0_valid; // @[extracted_function_conv.scala 143:31]
  wire [31:0] binaryOp_mul518_io_Out_0_bits_data; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_io_LeftIO_ready; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_io_LeftIO_valid; // @[extracted_function_conv.scala 143:31]
  wire [31:0] binaryOp_mul518_io_LeftIO_bits_data; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_io_RightIO_ready; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_mul518_io_RightIO_valid; // @[extracted_function_conv.scala 143:31]
  wire [31:0] binaryOp_mul518_io_RightIO_bits_data; // @[extracted_function_conv.scala 143:31]
  wire  binaryOp_sub619_clock; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_reset; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_io_enable_ready; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_io_enable_valid; // @[extracted_function_conv.scala 146:31]
  wire [4:0] binaryOp_sub619_io_enable_bits_taskID; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_io_enable_bits_control; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_io_Out_0_ready; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_io_Out_0_valid; // @[extracted_function_conv.scala 146:31]
  wire [31:0] binaryOp_sub619_io_Out_0_bits_data; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_io_LeftIO_ready; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_io_LeftIO_valid; // @[extracted_function_conv.scala 146:31]
  wire [31:0] binaryOp_sub619_io_LeftIO_bits_data; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_io_RightIO_ready; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_sub619_io_RightIO_valid; // @[extracted_function_conv.scala 146:31]
  wire [31:0] binaryOp_sub619_io_RightIO_bits_data; // @[extracted_function_conv.scala 146:31]
  wire  binaryOp_mul720_clock; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_reset; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_io_enable_ready; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_io_enable_valid; // @[extracted_function_conv.scala 149:31]
  wire [4:0] binaryOp_mul720_io_enable_bits_taskID; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_io_enable_bits_control; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_io_Out_0_ready; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_io_Out_0_valid; // @[extracted_function_conv.scala 149:31]
  wire [31:0] binaryOp_mul720_io_Out_0_bits_data; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_io_LeftIO_ready; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_io_LeftIO_valid; // @[extracted_function_conv.scala 149:31]
  wire [31:0] binaryOp_mul720_io_LeftIO_bits_data; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_io_RightIO_ready; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul720_io_RightIO_valid; // @[extracted_function_conv.scala 149:31]
  wire [31:0] binaryOp_mul720_io_RightIO_bits_data; // @[extracted_function_conv.scala 149:31]
  wire  binaryOp_mul821_clock; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_reset; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_io_enable_ready; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_io_enable_valid; // @[extracted_function_conv.scala 152:31]
  wire [4:0] binaryOp_mul821_io_enable_bits_taskID; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_io_enable_bits_control; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_io_Out_0_ready; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_io_Out_0_valid; // @[extracted_function_conv.scala 152:31]
  wire [31:0] binaryOp_mul821_io_Out_0_bits_data; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_io_LeftIO_ready; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_io_LeftIO_valid; // @[extracted_function_conv.scala 152:31]
  wire [31:0] binaryOp_mul821_io_LeftIO_bits_data; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_io_RightIO_ready; // @[extracted_function_conv.scala 152:31]
  wire  binaryOp_mul821_io_RightIO_valid; // @[extracted_function_conv.scala 152:31]
  wire  br_22_clock; // @[extracted_function_conv.scala 155:21]
  wire  br_22_reset; // @[extracted_function_conv.scala 155:21]
  wire  br_22_io_enable_ready; // @[extracted_function_conv.scala 155:21]
  wire  br_22_io_enable_valid; // @[extracted_function_conv.scala 155:21]
  wire [4:0] br_22_io_enable_bits_taskID; // @[extracted_function_conv.scala 155:21]
  wire  br_22_io_enable_bits_control; // @[extracted_function_conv.scala 155:21]
  wire  br_22_io_Out_0_ready; // @[extracted_function_conv.scala 155:21]
  wire  br_22_io_Out_0_valid; // @[extracted_function_conv.scala 155:21]
  wire [4:0] br_22_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 155:21]
  wire  br_22_io_Out_0_bits_control; // @[extracted_function_conv.scala 155:21]
  wire  binaryOp_inc12023_clock; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_reset; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_enable_ready; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_enable_valid; // @[extracted_function_conv.scala 158:33]
  wire [4:0] binaryOp_inc12023_io_enable_bits_taskID; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_enable_bits_control; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_Out_0_ready; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_Out_0_valid; // @[extracted_function_conv.scala 158:33]
  wire [4:0] binaryOp_inc12023_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 158:33]
  wire [31:0] binaryOp_inc12023_io_Out_0_bits_data; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_Out_1_ready; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_Out_1_valid; // @[extracted_function_conv.scala 158:33]
  wire [31:0] binaryOp_inc12023_io_Out_1_bits_data; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_LeftIO_ready; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_LeftIO_valid; // @[extracted_function_conv.scala 158:33]
  wire [31:0] binaryOp_inc12023_io_LeftIO_bits_data; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_RightIO_ready; // @[extracted_function_conv.scala 158:33]
  wire  binaryOp_inc12023_io_RightIO_valid; // @[extracted_function_conv.scala 158:33]
  wire  icmp_exitcond31424_clock; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_reset; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_io_enable_ready; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_io_enable_valid; // @[extracted_function_conv.scala 161:34]
  wire [4:0] icmp_exitcond31424_io_enable_bits_taskID; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_io_enable_bits_control; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_io_Out_0_ready; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_io_Out_0_valid; // @[extracted_function_conv.scala 161:34]
  wire [4:0] icmp_exitcond31424_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 161:34]
  wire [31:0] icmp_exitcond31424_io_Out_0_bits_data; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_io_LeftIO_ready; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_io_LeftIO_valid; // @[extracted_function_conv.scala 161:34]
  wire [31:0] icmp_exitcond31424_io_LeftIO_bits_data; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_io_RightIO_ready; // @[extracted_function_conv.scala 161:34]
  wire  icmp_exitcond31424_io_RightIO_valid; // @[extracted_function_conv.scala 161:34]
  wire  br_25_clock; // @[extracted_function_conv.scala 164:21]
  wire  br_25_reset; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_enable_ready; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_enable_valid; // @[extracted_function_conv.scala 164:21]
  wire [4:0] br_25_io_enable_bits_taskID; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_enable_bits_control; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_CmpIO_ready; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_CmpIO_valid; // @[extracted_function_conv.scala 164:21]
  wire [4:0] br_25_io_CmpIO_bits_taskID; // @[extracted_function_conv.scala 164:21]
  wire [31:0] br_25_io_CmpIO_bits_data; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_TrueOutput_0_ready; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_TrueOutput_0_valid; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_TrueOutput_0_bits_control; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_FalseOutput_0_ready; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_FalseOutput_0_valid; // @[extracted_function_conv.scala 164:21]
  wire [4:0] br_25_io_FalseOutput_0_bits_taskID; // @[extracted_function_conv.scala 164:21]
  wire  br_25_io_FalseOutput_0_bits_control; // @[extracted_function_conv.scala 164:21]
  wire  phi_conv_s1_x_031226_clock; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_reset; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_enable_ready; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_enable_valid; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_enable_bits_control; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_InData_0_ready; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_InData_0_valid; // @[extracted_function_conv.scala 167:36]
  wire [4:0] phi_conv_s1_x_031226_io_InData_0_bits_taskID; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_InData_1_ready; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_InData_1_valid; // @[extracted_function_conv.scala 167:36]
  wire [4:0] phi_conv_s1_x_031226_io_InData_1_bits_taskID; // @[extracted_function_conv.scala 167:36]
  wire [31:0] phi_conv_s1_x_031226_io_InData_1_bits_data; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Mask_ready; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Mask_valid; // @[extracted_function_conv.scala 167:36]
  wire [1:0] phi_conv_s1_x_031226_io_Mask_bits; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Out_0_ready; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Out_0_valid; // @[extracted_function_conv.scala 167:36]
  wire [31:0] phi_conv_s1_x_031226_io_Out_0_bits_data; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Out_1_ready; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Out_1_valid; // @[extracted_function_conv.scala 167:36]
  wire [31:0] phi_conv_s1_x_031226_io_Out_1_bits_data; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Out_2_ready; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Out_2_valid; // @[extracted_function_conv.scala 167:36]
  wire [31:0] phi_conv_s1_x_031226_io_Out_2_bits_data; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Out_3_ready; // @[extracted_function_conv.scala 167:36]
  wire  phi_conv_s1_x_031226_io_Out_3_valid; // @[extracted_function_conv.scala 167:36]
  wire [31:0] phi_conv_s1_x_031226_io_Out_3_bits_data; // @[extracted_function_conv.scala 167:36]
  wire  binaryOp_add1327_clock; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_reset; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_io_enable_ready; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_io_enable_valid; // @[extracted_function_conv.scala 170:32]
  wire [4:0] binaryOp_add1327_io_enable_bits_taskID; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_io_enable_bits_control; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_io_Out_0_ready; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_io_Out_0_valid; // @[extracted_function_conv.scala 170:32]
  wire [31:0] binaryOp_add1327_io_Out_0_bits_data; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_io_LeftIO_ready; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_io_LeftIO_valid; // @[extracted_function_conv.scala 170:32]
  wire [31:0] binaryOp_add1327_io_LeftIO_bits_data; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_io_RightIO_ready; // @[extracted_function_conv.scala 170:32]
  wire  binaryOp_add1327_io_RightIO_valid; // @[extracted_function_conv.scala 170:32]
  wire [31:0] binaryOp_add1327_io_RightIO_bits_data; // @[extracted_function_conv.scala 170:32]
  wire  Gep_arrayidx28_clock; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_reset; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_enable_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_enable_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_enable_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_enable_bits_control; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_0_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_0_valid; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_0_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_1_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_1_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_1_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_2_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_2_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_2_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_3_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_3_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_3_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_4_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_4_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_4_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_5_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_5_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_5_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_5_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_6_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_6_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_6_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_6_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_7_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_7_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_7_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_7_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_8_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_8_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_8_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_8_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_9_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_Out_9_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_Out_9_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_Out_9_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_baseAddress_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_baseAddress_valid; // @[extracted_function_conv.scala 173:30]
  wire [4:0] Gep_arrayidx28_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_baseAddress_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_idx_0_ready; // @[extracted_function_conv.scala 173:30]
  wire  Gep_arrayidx28_io_idx_0_valid; // @[extracted_function_conv.scala 173:30]
  wire [31:0] Gep_arrayidx28_io_idx_0_bits_data; // @[extracted_function_conv.scala 173:30]
  wire  ld_29_clock; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_reset; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_enable_ready; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_enable_valid; // @[extracted_function_conv.scala 176:21]
  wire [4:0] ld_29_io_enable_bits_taskID; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_enable_bits_control; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_Out_0_ready; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_Out_0_valid; // @[extracted_function_conv.scala 176:21]
  wire [31:0] ld_29_io_Out_0_bits_data; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_GepAddr_ready; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_GepAddr_valid; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 176:21]
  wire [4:0] ld_29_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 176:21]
  wire [31:0] ld_29_io_GepAddr_bits_data; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_memReq_ready; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_memReq_valid; // @[extracted_function_conv.scala 176:21]
  wire [31:0] ld_29_io_memReq_bits_address; // @[extracted_function_conv.scala 176:21]
  wire [4:0] ld_29_io_memReq_bits_taskID; // @[extracted_function_conv.scala 176:21]
  wire  ld_29_io_memResp_valid; // @[extracted_function_conv.scala 176:21]
  wire [31:0] ld_29_io_memResp_data; // @[extracted_function_conv.scala 176:21]
  wire  ld_30_clock; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_reset; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_enable_ready; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_enable_valid; // @[extracted_function_conv.scala 179:21]
  wire [4:0] ld_30_io_enable_bits_taskID; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_enable_bits_control; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_Out_0_ready; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_Out_0_valid; // @[extracted_function_conv.scala 179:21]
  wire [31:0] ld_30_io_Out_0_bits_data; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_GepAddr_ready; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_GepAddr_valid; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 179:21]
  wire [4:0] ld_30_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 179:21]
  wire [31:0] ld_30_io_GepAddr_bits_data; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_memReq_ready; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_memReq_valid; // @[extracted_function_conv.scala 179:21]
  wire [31:0] ld_30_io_memReq_bits_address; // @[extracted_function_conv.scala 179:21]
  wire [4:0] ld_30_io_memReq_bits_taskID; // @[extracted_function_conv.scala 179:21]
  wire  ld_30_io_memResp_valid; // @[extracted_function_conv.scala 179:21]
  wire [31:0] ld_30_io_memResp_data; // @[extracted_function_conv.scala 179:21]
  wire  binaryOp_add1531_clock; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_reset; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_io_enable_ready; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_io_enable_valid; // @[extracted_function_conv.scala 182:32]
  wire [4:0] binaryOp_add1531_io_enable_bits_taskID; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_io_enable_bits_control; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_io_Out_0_ready; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_io_Out_0_valid; // @[extracted_function_conv.scala 182:32]
  wire [31:0] binaryOp_add1531_io_Out_0_bits_data; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_io_LeftIO_ready; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_io_LeftIO_valid; // @[extracted_function_conv.scala 182:32]
  wire [31:0] binaryOp_add1531_io_LeftIO_bits_data; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_io_RightIO_ready; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_add1531_io_RightIO_valid; // @[extracted_function_conv.scala 182:32]
  wire [31:0] binaryOp_add1531_io_RightIO_bits_data; // @[extracted_function_conv.scala 182:32]
  wire  binaryOp_mul1632_clock; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_reset; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_io_enable_ready; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_io_enable_valid; // @[extracted_function_conv.scala 185:32]
  wire [4:0] binaryOp_mul1632_io_enable_bits_taskID; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_io_enable_bits_control; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_io_Out_0_ready; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_io_Out_0_valid; // @[extracted_function_conv.scala 185:32]
  wire [31:0] binaryOp_mul1632_io_Out_0_bits_data; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_io_LeftIO_ready; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_io_LeftIO_valid; // @[extracted_function_conv.scala 185:32]
  wire [31:0] binaryOp_mul1632_io_LeftIO_bits_data; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_io_RightIO_ready; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_mul1632_io_RightIO_valid; // @[extracted_function_conv.scala 185:32]
  wire  binaryOp_sub1733_clock; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_reset; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_enable_ready; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_enable_valid; // @[extracted_function_conv.scala 188:32]
  wire [4:0] binaryOp_sub1733_io_enable_bits_taskID; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_enable_bits_control; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_Out_0_ready; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_Out_0_valid; // @[extracted_function_conv.scala 188:32]
  wire [31:0] binaryOp_sub1733_io_Out_0_bits_data; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_Out_1_ready; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_Out_1_valid; // @[extracted_function_conv.scala 188:32]
  wire [31:0] binaryOp_sub1733_io_Out_1_bits_data; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_Out_2_ready; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_Out_2_valid; // @[extracted_function_conv.scala 188:32]
  wire [31:0] binaryOp_sub1733_io_Out_2_bits_data; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_LeftIO_ready; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_LeftIO_valid; // @[extracted_function_conv.scala 188:32]
  wire [31:0] binaryOp_sub1733_io_LeftIO_bits_data; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_RightIO_ready; // @[extracted_function_conv.scala 188:32]
  wire  binaryOp_sub1733_io_RightIO_valid; // @[extracted_function_conv.scala 188:32]
  wire [31:0] binaryOp_sub1733_io_RightIO_bits_data; // @[extracted_function_conv.scala 188:32]
  wire  Gep_arrayidx1834_clock; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_reset; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_enable_ready; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_enable_valid; // @[extracted_function_conv.scala 191:32]
  wire [4:0] Gep_arrayidx1834_io_enable_bits_taskID; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_enable_bits_control; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_Out_0_ready; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_Out_0_valid; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 191:32]
  wire [4:0] Gep_arrayidx1834_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 191:32]
  wire [31:0] Gep_arrayidx1834_io_Out_0_bits_data; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_baseAddress_ready; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_baseAddress_valid; // @[extracted_function_conv.scala 191:32]
  wire [4:0] Gep_arrayidx1834_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 191:32]
  wire [31:0] Gep_arrayidx1834_io_baseAddress_bits_data; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_idx_0_ready; // @[extracted_function_conv.scala 191:32]
  wire  Gep_arrayidx1834_io_idx_0_valid; // @[extracted_function_conv.scala 191:32]
  wire [31:0] Gep_arrayidx1834_io_idx_0_bits_data; // @[extracted_function_conv.scala 191:32]
  wire  ld_35_clock; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_reset; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_enable_ready; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_enable_valid; // @[extracted_function_conv.scala 194:21]
  wire [4:0] ld_35_io_enable_bits_taskID; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_enable_bits_control; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_Out_0_ready; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_Out_0_valid; // @[extracted_function_conv.scala 194:21]
  wire [31:0] ld_35_io_Out_0_bits_data; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_GepAddr_ready; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_GepAddr_valid; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 194:21]
  wire [4:0] ld_35_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 194:21]
  wire [31:0] ld_35_io_GepAddr_bits_data; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_memReq_ready; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_memReq_valid; // @[extracted_function_conv.scala 194:21]
  wire [31:0] ld_35_io_memReq_bits_address; // @[extracted_function_conv.scala 194:21]
  wire [4:0] ld_35_io_memReq_bits_taskID; // @[extracted_function_conv.scala 194:21]
  wire  ld_35_io_memResp_valid; // @[extracted_function_conv.scala 194:21]
  wire [31:0] ld_35_io_memResp_data; // @[extracted_function_conv.scala 194:21]
  wire  sextconv1936_clock; // @[extracted_function_conv.scala 197:28]
  wire  sextconv1936_reset; // @[extracted_function_conv.scala 197:28]
  wire  sextconv1936_io_Input_ready; // @[extracted_function_conv.scala 197:28]
  wire  sextconv1936_io_Input_valid; // @[extracted_function_conv.scala 197:28]
  wire [31:0] sextconv1936_io_Input_bits_data; // @[extracted_function_conv.scala 197:28]
  wire  sextconv1936_io_enable_ready; // @[extracted_function_conv.scala 197:28]
  wire  sextconv1936_io_enable_valid; // @[extracted_function_conv.scala 197:28]
  wire [4:0] sextconv1936_io_enable_bits_taskID; // @[extracted_function_conv.scala 197:28]
  wire  sextconv1936_io_Out_0_ready; // @[extracted_function_conv.scala 197:28]
  wire  sextconv1936_io_Out_0_valid; // @[extracted_function_conv.scala 197:28]
  wire [31:0] sextconv1936_io_Out_0_bits_data; // @[extracted_function_conv.scala 197:28]
  wire  binaryOp_mul2037_clock; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_reset; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_io_enable_ready; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_io_enable_valid; // @[extracted_function_conv.scala 200:32]
  wire [4:0] binaryOp_mul2037_io_enable_bits_taskID; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_io_enable_bits_control; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_io_Out_0_ready; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_io_Out_0_valid; // @[extracted_function_conv.scala 200:32]
  wire [31:0] binaryOp_mul2037_io_Out_0_bits_data; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_io_LeftIO_ready; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_io_LeftIO_valid; // @[extracted_function_conv.scala 200:32]
  wire [31:0] binaryOp_mul2037_io_LeftIO_bits_data; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_io_RightIO_ready; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_mul2037_io_RightIO_valid; // @[extracted_function_conv.scala 200:32]
  wire [31:0] binaryOp_mul2037_io_RightIO_bits_data; // @[extracted_function_conv.scala 200:32]
  wire  binaryOp_add2138_clock; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_reset; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_enable_ready; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_enable_valid; // @[extracted_function_conv.scala 203:32]
  wire [4:0] binaryOp_add2138_io_enable_bits_taskID; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_enable_bits_control; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_Out_0_ready; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_Out_0_valid; // @[extracted_function_conv.scala 203:32]
  wire [4:0] binaryOp_add2138_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 203:32]
  wire [31:0] binaryOp_add2138_io_Out_0_bits_data; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_Out_1_ready; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_Out_1_valid; // @[extracted_function_conv.scala 203:32]
  wire [31:0] binaryOp_add2138_io_Out_1_bits_data; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_LeftIO_ready; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_LeftIO_valid; // @[extracted_function_conv.scala 203:32]
  wire [31:0] binaryOp_add2138_io_LeftIO_bits_data; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_RightIO_ready; // @[extracted_function_conv.scala 203:32]
  wire  binaryOp_add2138_io_RightIO_valid; // @[extracted_function_conv.scala 203:32]
  wire [31:0] binaryOp_add2138_io_RightIO_bits_data; // @[extracted_function_conv.scala 203:32]
  wire  st_39_clock; // @[extracted_function_conv.scala 206:21]
  wire  st_39_reset; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_enable_ready; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_enable_valid; // @[extracted_function_conv.scala 206:21]
  wire [4:0] st_39_io_enable_bits_taskID; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_enable_bits_control; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_GepAddr_ready; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_GepAddr_valid; // @[extracted_function_conv.scala 206:21]
  wire [4:0] st_39_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 206:21]
  wire [31:0] st_39_io_GepAddr_bits_data; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_inData_ready; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_inData_valid; // @[extracted_function_conv.scala 206:21]
  wire [4:0] st_39_io_inData_bits_taskID; // @[extracted_function_conv.scala 206:21]
  wire [31:0] st_39_io_inData_bits_data; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_memReq_ready; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_memReq_valid; // @[extracted_function_conv.scala 206:21]
  wire [21:0] st_39_io_memReq_bits_address; // @[extracted_function_conv.scala 206:21]
  wire [31:0] st_39_io_memReq_bits_data; // @[extracted_function_conv.scala 206:21]
  wire [4:0] st_39_io_memReq_bits_taskID; // @[extracted_function_conv.scala 206:21]
  wire  st_39_io_memResp_valid; // @[extracted_function_conv.scala 206:21]
  wire  ld_40_clock; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_reset; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_enable_ready; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_enable_valid; // @[extracted_function_conv.scala 209:21]
  wire [4:0] ld_40_io_enable_bits_taskID; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_enable_bits_control; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_Out_0_ready; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_Out_0_valid; // @[extracted_function_conv.scala 209:21]
  wire [31:0] ld_40_io_Out_0_bits_data; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_GepAddr_ready; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_GepAddr_valid; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 209:21]
  wire [4:0] ld_40_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 209:21]
  wire [31:0] ld_40_io_GepAddr_bits_data; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_memReq_ready; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_memReq_valid; // @[extracted_function_conv.scala 209:21]
  wire [31:0] ld_40_io_memReq_bits_address; // @[extracted_function_conv.scala 209:21]
  wire [4:0] ld_40_io_memReq_bits_taskID; // @[extracted_function_conv.scala 209:21]
  wire  ld_40_io_memResp_valid; // @[extracted_function_conv.scala 209:21]
  wire [31:0] ld_40_io_memResp_data; // @[extracted_function_conv.scala 209:21]
  wire  binaryOp_add2941_clock; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_reset; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_io_enable_ready; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_io_enable_valid; // @[extracted_function_conv.scala 212:32]
  wire [4:0] binaryOp_add2941_io_enable_bits_taskID; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_io_enable_bits_control; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_io_Out_0_ready; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_io_Out_0_valid; // @[extracted_function_conv.scala 212:32]
  wire [31:0] binaryOp_add2941_io_Out_0_bits_data; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_io_LeftIO_ready; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_io_LeftIO_valid; // @[extracted_function_conv.scala 212:32]
  wire [31:0] binaryOp_add2941_io_LeftIO_bits_data; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_io_RightIO_ready; // @[extracted_function_conv.scala 212:32]
  wire  binaryOp_add2941_io_RightIO_valid; // @[extracted_function_conv.scala 212:32]
  wire  Gep_arrayidx3042_clock; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_reset; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_enable_ready; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_enable_valid; // @[extracted_function_conv.scala 215:32]
  wire [4:0] Gep_arrayidx3042_io_enable_bits_taskID; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_enable_bits_control; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_Out_0_ready; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_Out_0_valid; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 215:32]
  wire [4:0] Gep_arrayidx3042_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 215:32]
  wire [31:0] Gep_arrayidx3042_io_Out_0_bits_data; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_baseAddress_ready; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_baseAddress_valid; // @[extracted_function_conv.scala 215:32]
  wire [4:0] Gep_arrayidx3042_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 215:32]
  wire [31:0] Gep_arrayidx3042_io_baseAddress_bits_data; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_idx_0_ready; // @[extracted_function_conv.scala 215:32]
  wire  Gep_arrayidx3042_io_idx_0_valid; // @[extracted_function_conv.scala 215:32]
  wire [31:0] Gep_arrayidx3042_io_idx_0_bits_data; // @[extracted_function_conv.scala 215:32]
  wire  ld_43_clock; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_reset; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_enable_ready; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_enable_valid; // @[extracted_function_conv.scala 218:21]
  wire [4:0] ld_43_io_enable_bits_taskID; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_enable_bits_control; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_Out_0_ready; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_Out_0_valid; // @[extracted_function_conv.scala 218:21]
  wire [31:0] ld_43_io_Out_0_bits_data; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_GepAddr_ready; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_GepAddr_valid; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 218:21]
  wire [4:0] ld_43_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 218:21]
  wire [31:0] ld_43_io_GepAddr_bits_data; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_memReq_ready; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_memReq_valid; // @[extracted_function_conv.scala 218:21]
  wire [31:0] ld_43_io_memReq_bits_address; // @[extracted_function_conv.scala 218:21]
  wire [4:0] ld_43_io_memReq_bits_taskID; // @[extracted_function_conv.scala 218:21]
  wire  ld_43_io_memResp_valid; // @[extracted_function_conv.scala 218:21]
  wire [31:0] ld_43_io_memResp_data; // @[extracted_function_conv.scala 218:21]
  wire  sextconv3244_clock; // @[extracted_function_conv.scala 221:28]
  wire  sextconv3244_reset; // @[extracted_function_conv.scala 221:28]
  wire  sextconv3244_io_Input_ready; // @[extracted_function_conv.scala 221:28]
  wire  sextconv3244_io_Input_valid; // @[extracted_function_conv.scala 221:28]
  wire [31:0] sextconv3244_io_Input_bits_data; // @[extracted_function_conv.scala 221:28]
  wire  sextconv3244_io_enable_ready; // @[extracted_function_conv.scala 221:28]
  wire  sextconv3244_io_enable_valid; // @[extracted_function_conv.scala 221:28]
  wire [4:0] sextconv3244_io_enable_bits_taskID; // @[extracted_function_conv.scala 221:28]
  wire  sextconv3244_io_Out_0_ready; // @[extracted_function_conv.scala 221:28]
  wire  sextconv3244_io_Out_0_valid; // @[extracted_function_conv.scala 221:28]
  wire [31:0] sextconv3244_io_Out_0_bits_data; // @[extracted_function_conv.scala 221:28]
  wire  binaryOp_mul3345_clock; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_reset; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_io_enable_ready; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_io_enable_valid; // @[extracted_function_conv.scala 224:32]
  wire [4:0] binaryOp_mul3345_io_enable_bits_taskID; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_io_enable_bits_control; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_io_Out_0_ready; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_io_Out_0_valid; // @[extracted_function_conv.scala 224:32]
  wire [31:0] binaryOp_mul3345_io_Out_0_bits_data; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_io_LeftIO_ready; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_io_LeftIO_valid; // @[extracted_function_conv.scala 224:32]
  wire [31:0] binaryOp_mul3345_io_LeftIO_bits_data; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_io_RightIO_ready; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_mul3345_io_RightIO_valid; // @[extracted_function_conv.scala 224:32]
  wire [31:0] binaryOp_mul3345_io_RightIO_bits_data; // @[extracted_function_conv.scala 224:32]
  wire  binaryOp_add3446_clock; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_reset; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_enable_ready; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_enable_valid; // @[extracted_function_conv.scala 227:32]
  wire [4:0] binaryOp_add3446_io_enable_bits_taskID; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_enable_bits_control; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_Out_0_ready; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_Out_0_valid; // @[extracted_function_conv.scala 227:32]
  wire [4:0] binaryOp_add3446_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 227:32]
  wire [31:0] binaryOp_add3446_io_Out_0_bits_data; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_Out_1_ready; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_Out_1_valid; // @[extracted_function_conv.scala 227:32]
  wire [31:0] binaryOp_add3446_io_Out_1_bits_data; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_LeftIO_ready; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_LeftIO_valid; // @[extracted_function_conv.scala 227:32]
  wire [31:0] binaryOp_add3446_io_LeftIO_bits_data; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_RightIO_ready; // @[extracted_function_conv.scala 227:32]
  wire  binaryOp_add3446_io_RightIO_valid; // @[extracted_function_conv.scala 227:32]
  wire [31:0] binaryOp_add3446_io_RightIO_bits_data; // @[extracted_function_conv.scala 227:32]
  wire  st_47_clock; // @[extracted_function_conv.scala 230:21]
  wire  st_47_reset; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_enable_ready; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_enable_valid; // @[extracted_function_conv.scala 230:21]
  wire [4:0] st_47_io_enable_bits_taskID; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_enable_bits_control; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_GepAddr_ready; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_GepAddr_valid; // @[extracted_function_conv.scala 230:21]
  wire [4:0] st_47_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 230:21]
  wire [31:0] st_47_io_GepAddr_bits_data; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_inData_ready; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_inData_valid; // @[extracted_function_conv.scala 230:21]
  wire [4:0] st_47_io_inData_bits_taskID; // @[extracted_function_conv.scala 230:21]
  wire [31:0] st_47_io_inData_bits_data; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_memReq_ready; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_memReq_valid; // @[extracted_function_conv.scala 230:21]
  wire [21:0] st_47_io_memReq_bits_address; // @[extracted_function_conv.scala 230:21]
  wire [31:0] st_47_io_memReq_bits_data; // @[extracted_function_conv.scala 230:21]
  wire [4:0] st_47_io_memReq_bits_taskID; // @[extracted_function_conv.scala 230:21]
  wire  st_47_io_memResp_valid; // @[extracted_function_conv.scala 230:21]
  wire  ld_48_clock; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_reset; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_enable_ready; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_enable_valid; // @[extracted_function_conv.scala 233:21]
  wire [4:0] ld_48_io_enable_bits_taskID; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_enable_bits_control; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_Out_0_ready; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_Out_0_valid; // @[extracted_function_conv.scala 233:21]
  wire [31:0] ld_48_io_Out_0_bits_data; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_GepAddr_ready; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_GepAddr_valid; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 233:21]
  wire [4:0] ld_48_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 233:21]
  wire [31:0] ld_48_io_GepAddr_bits_data; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_memReq_ready; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_memReq_valid; // @[extracted_function_conv.scala 233:21]
  wire [31:0] ld_48_io_memReq_bits_address; // @[extracted_function_conv.scala 233:21]
  wire [4:0] ld_48_io_memReq_bits_taskID; // @[extracted_function_conv.scala 233:21]
  wire  ld_48_io_memResp_valid; // @[extracted_function_conv.scala 233:21]
  wire [31:0] ld_48_io_memResp_data; // @[extracted_function_conv.scala 233:21]
  wire  binaryOp_add4249_clock; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_reset; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_io_enable_ready; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_io_enable_valid; // @[extracted_function_conv.scala 236:32]
  wire [4:0] binaryOp_add4249_io_enable_bits_taskID; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_io_enable_bits_control; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_io_Out_0_ready; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_io_Out_0_valid; // @[extracted_function_conv.scala 236:32]
  wire [31:0] binaryOp_add4249_io_Out_0_bits_data; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_io_LeftIO_ready; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_io_LeftIO_valid; // @[extracted_function_conv.scala 236:32]
  wire [31:0] binaryOp_add4249_io_LeftIO_bits_data; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_io_RightIO_ready; // @[extracted_function_conv.scala 236:32]
  wire  binaryOp_add4249_io_RightIO_valid; // @[extracted_function_conv.scala 236:32]
  wire  Gep_arrayidx4350_clock; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_reset; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_enable_ready; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_enable_valid; // @[extracted_function_conv.scala 239:32]
  wire [4:0] Gep_arrayidx4350_io_enable_bits_taskID; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_enable_bits_control; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_Out_0_ready; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_Out_0_valid; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 239:32]
  wire [4:0] Gep_arrayidx4350_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 239:32]
  wire [31:0] Gep_arrayidx4350_io_Out_0_bits_data; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_baseAddress_ready; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_baseAddress_valid; // @[extracted_function_conv.scala 239:32]
  wire [4:0] Gep_arrayidx4350_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 239:32]
  wire [31:0] Gep_arrayidx4350_io_baseAddress_bits_data; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_idx_0_ready; // @[extracted_function_conv.scala 239:32]
  wire  Gep_arrayidx4350_io_idx_0_valid; // @[extracted_function_conv.scala 239:32]
  wire [31:0] Gep_arrayidx4350_io_idx_0_bits_data; // @[extracted_function_conv.scala 239:32]
  wire  ld_51_clock; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_reset; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_enable_ready; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_enable_valid; // @[extracted_function_conv.scala 242:21]
  wire [4:0] ld_51_io_enable_bits_taskID; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_enable_bits_control; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_Out_0_ready; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_Out_0_valid; // @[extracted_function_conv.scala 242:21]
  wire [31:0] ld_51_io_Out_0_bits_data; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_GepAddr_ready; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_GepAddr_valid; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 242:21]
  wire [4:0] ld_51_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 242:21]
  wire [31:0] ld_51_io_GepAddr_bits_data; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_memReq_ready; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_memReq_valid; // @[extracted_function_conv.scala 242:21]
  wire [31:0] ld_51_io_memReq_bits_address; // @[extracted_function_conv.scala 242:21]
  wire [4:0] ld_51_io_memReq_bits_taskID; // @[extracted_function_conv.scala 242:21]
  wire  ld_51_io_memResp_valid; // @[extracted_function_conv.scala 242:21]
  wire [31:0] ld_51_io_memResp_data; // @[extracted_function_conv.scala 242:21]
  wire  sextconv4552_clock; // @[extracted_function_conv.scala 245:28]
  wire  sextconv4552_reset; // @[extracted_function_conv.scala 245:28]
  wire  sextconv4552_io_Input_ready; // @[extracted_function_conv.scala 245:28]
  wire  sextconv4552_io_Input_valid; // @[extracted_function_conv.scala 245:28]
  wire [31:0] sextconv4552_io_Input_bits_data; // @[extracted_function_conv.scala 245:28]
  wire  sextconv4552_io_enable_ready; // @[extracted_function_conv.scala 245:28]
  wire  sextconv4552_io_enable_valid; // @[extracted_function_conv.scala 245:28]
  wire [4:0] sextconv4552_io_enable_bits_taskID; // @[extracted_function_conv.scala 245:28]
  wire  sextconv4552_io_Out_0_ready; // @[extracted_function_conv.scala 245:28]
  wire  sextconv4552_io_Out_0_valid; // @[extracted_function_conv.scala 245:28]
  wire [31:0] sextconv4552_io_Out_0_bits_data; // @[extracted_function_conv.scala 245:28]
  wire  binaryOp_mul4653_clock; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_reset; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_io_enable_ready; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_io_enable_valid; // @[extracted_function_conv.scala 248:32]
  wire [4:0] binaryOp_mul4653_io_enable_bits_taskID; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_io_enable_bits_control; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_io_Out_0_ready; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_io_Out_0_valid; // @[extracted_function_conv.scala 248:32]
  wire [31:0] binaryOp_mul4653_io_Out_0_bits_data; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_io_LeftIO_ready; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_io_LeftIO_valid; // @[extracted_function_conv.scala 248:32]
  wire [31:0] binaryOp_mul4653_io_LeftIO_bits_data; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_io_RightIO_ready; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_mul4653_io_RightIO_valid; // @[extracted_function_conv.scala 248:32]
  wire [31:0] binaryOp_mul4653_io_RightIO_bits_data; // @[extracted_function_conv.scala 248:32]
  wire  binaryOp_add4754_clock; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_reset; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_enable_ready; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_enable_valid; // @[extracted_function_conv.scala 251:32]
  wire [4:0] binaryOp_add4754_io_enable_bits_taskID; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_enable_bits_control; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_Out_0_ready; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_Out_0_valid; // @[extracted_function_conv.scala 251:32]
  wire [4:0] binaryOp_add4754_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 251:32]
  wire [31:0] binaryOp_add4754_io_Out_0_bits_data; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_Out_1_ready; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_Out_1_valid; // @[extracted_function_conv.scala 251:32]
  wire [31:0] binaryOp_add4754_io_Out_1_bits_data; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_LeftIO_ready; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_LeftIO_valid; // @[extracted_function_conv.scala 251:32]
  wire [31:0] binaryOp_add4754_io_LeftIO_bits_data; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_RightIO_ready; // @[extracted_function_conv.scala 251:32]
  wire  binaryOp_add4754_io_RightIO_valid; // @[extracted_function_conv.scala 251:32]
  wire [31:0] binaryOp_add4754_io_RightIO_bits_data; // @[extracted_function_conv.scala 251:32]
  wire  st_55_clock; // @[extracted_function_conv.scala 254:21]
  wire  st_55_reset; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_enable_ready; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_enable_valid; // @[extracted_function_conv.scala 254:21]
  wire [4:0] st_55_io_enable_bits_taskID; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_enable_bits_control; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_GepAddr_ready; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_GepAddr_valid; // @[extracted_function_conv.scala 254:21]
  wire [4:0] st_55_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 254:21]
  wire [31:0] st_55_io_GepAddr_bits_data; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_inData_ready; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_inData_valid; // @[extracted_function_conv.scala 254:21]
  wire [4:0] st_55_io_inData_bits_taskID; // @[extracted_function_conv.scala 254:21]
  wire [31:0] st_55_io_inData_bits_data; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_memReq_ready; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_memReq_valid; // @[extracted_function_conv.scala 254:21]
  wire [21:0] st_55_io_memReq_bits_address; // @[extracted_function_conv.scala 254:21]
  wire [31:0] st_55_io_memReq_bits_data; // @[extracted_function_conv.scala 254:21]
  wire [4:0] st_55_io_memReq_bits_taskID; // @[extracted_function_conv.scala 254:21]
  wire  st_55_io_memResp_valid; // @[extracted_function_conv.scala 254:21]
  wire  ld_56_clock; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_reset; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_enable_ready; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_enable_valid; // @[extracted_function_conv.scala 257:21]
  wire [4:0] ld_56_io_enable_bits_taskID; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_enable_bits_control; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_Out_0_ready; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_Out_0_valid; // @[extracted_function_conv.scala 257:21]
  wire [31:0] ld_56_io_Out_0_bits_data; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_GepAddr_ready; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_GepAddr_valid; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 257:21]
  wire [4:0] ld_56_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 257:21]
  wire [31:0] ld_56_io_GepAddr_bits_data; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_memReq_ready; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_memReq_valid; // @[extracted_function_conv.scala 257:21]
  wire [31:0] ld_56_io_memReq_bits_address; // @[extracted_function_conv.scala 257:21]
  wire [4:0] ld_56_io_memReq_bits_taskID; // @[extracted_function_conv.scala 257:21]
  wire  ld_56_io_memResp_valid; // @[extracted_function_conv.scala 257:21]
  wire [31:0] ld_56_io_memResp_data; // @[extracted_function_conv.scala 257:21]
  wire  binaryOp_mul5257_clock; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_reset; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_enable_ready; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_enable_valid; // @[extracted_function_conv.scala 260:32]
  wire [4:0] binaryOp_mul5257_io_enable_bits_taskID; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_enable_bits_control; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_Out_0_ready; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_Out_0_valid; // @[extracted_function_conv.scala 260:32]
  wire [31:0] binaryOp_mul5257_io_Out_0_bits_data; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_Out_1_ready; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_Out_1_valid; // @[extracted_function_conv.scala 260:32]
  wire [31:0] binaryOp_mul5257_io_Out_1_bits_data; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_LeftIO_ready; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_LeftIO_valid; // @[extracted_function_conv.scala 260:32]
  wire [31:0] binaryOp_mul5257_io_LeftIO_bits_data; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_RightIO_ready; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_mul5257_io_RightIO_valid; // @[extracted_function_conv.scala 260:32]
  wire  binaryOp_add5358_clock; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_reset; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_enable_ready; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_enable_valid; // @[extracted_function_conv.scala 263:32]
  wire [4:0] binaryOp_add5358_io_enable_bits_taskID; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_enable_bits_control; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_Out_0_ready; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_Out_0_valid; // @[extracted_function_conv.scala 263:32]
  wire [31:0] binaryOp_add5358_io_Out_0_bits_data; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_Out_1_ready; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_Out_1_valid; // @[extracted_function_conv.scala 263:32]
  wire [31:0] binaryOp_add5358_io_Out_1_bits_data; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_Out_2_ready; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_Out_2_valid; // @[extracted_function_conv.scala 263:32]
  wire [31:0] binaryOp_add5358_io_Out_2_bits_data; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_LeftIO_ready; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_LeftIO_valid; // @[extracted_function_conv.scala 263:32]
  wire [31:0] binaryOp_add5358_io_LeftIO_bits_data; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_RightIO_ready; // @[extracted_function_conv.scala 263:32]
  wire  binaryOp_add5358_io_RightIO_valid; // @[extracted_function_conv.scala 263:32]
  wire [31:0] binaryOp_add5358_io_RightIO_bits_data; // @[extracted_function_conv.scala 263:32]
  wire  Gep_arrayidx5459_clock; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_reset; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_enable_ready; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_enable_valid; // @[extracted_function_conv.scala 266:32]
  wire [4:0] Gep_arrayidx5459_io_enable_bits_taskID; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_enable_bits_control; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_Out_0_ready; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_Out_0_valid; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 266:32]
  wire [4:0] Gep_arrayidx5459_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 266:32]
  wire [31:0] Gep_arrayidx5459_io_Out_0_bits_data; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_baseAddress_ready; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_baseAddress_valid; // @[extracted_function_conv.scala 266:32]
  wire [4:0] Gep_arrayidx5459_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 266:32]
  wire [31:0] Gep_arrayidx5459_io_baseAddress_bits_data; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_idx_0_ready; // @[extracted_function_conv.scala 266:32]
  wire  Gep_arrayidx5459_io_idx_0_valid; // @[extracted_function_conv.scala 266:32]
  wire [31:0] Gep_arrayidx5459_io_idx_0_bits_data; // @[extracted_function_conv.scala 266:32]
  wire  ld_60_clock; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_reset; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_enable_ready; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_enable_valid; // @[extracted_function_conv.scala 269:21]
  wire [4:0] ld_60_io_enable_bits_taskID; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_enable_bits_control; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_Out_0_ready; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_Out_0_valid; // @[extracted_function_conv.scala 269:21]
  wire [31:0] ld_60_io_Out_0_bits_data; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_GepAddr_ready; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_GepAddr_valid; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 269:21]
  wire [4:0] ld_60_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 269:21]
  wire [31:0] ld_60_io_GepAddr_bits_data; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_memReq_ready; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_memReq_valid; // @[extracted_function_conv.scala 269:21]
  wire [31:0] ld_60_io_memReq_bits_address; // @[extracted_function_conv.scala 269:21]
  wire [4:0] ld_60_io_memReq_bits_taskID; // @[extracted_function_conv.scala 269:21]
  wire  ld_60_io_memResp_valid; // @[extracted_function_conv.scala 269:21]
  wire [31:0] ld_60_io_memResp_data; // @[extracted_function_conv.scala 269:21]
  wire  sextconv5661_clock; // @[extracted_function_conv.scala 272:28]
  wire  sextconv5661_reset; // @[extracted_function_conv.scala 272:28]
  wire  sextconv5661_io_Input_ready; // @[extracted_function_conv.scala 272:28]
  wire  sextconv5661_io_Input_valid; // @[extracted_function_conv.scala 272:28]
  wire [31:0] sextconv5661_io_Input_bits_data; // @[extracted_function_conv.scala 272:28]
  wire  sextconv5661_io_enable_ready; // @[extracted_function_conv.scala 272:28]
  wire  sextconv5661_io_enable_valid; // @[extracted_function_conv.scala 272:28]
  wire [4:0] sextconv5661_io_enable_bits_taskID; // @[extracted_function_conv.scala 272:28]
  wire  sextconv5661_io_Out_0_ready; // @[extracted_function_conv.scala 272:28]
  wire  sextconv5661_io_Out_0_valid; // @[extracted_function_conv.scala 272:28]
  wire [31:0] sextconv5661_io_Out_0_bits_data; // @[extracted_function_conv.scala 272:28]
  wire  binaryOp_mul5762_clock; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_reset; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_io_enable_ready; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_io_enable_valid; // @[extracted_function_conv.scala 275:32]
  wire [4:0] binaryOp_mul5762_io_enable_bits_taskID; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_io_enable_bits_control; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_io_Out_0_ready; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_io_Out_0_valid; // @[extracted_function_conv.scala 275:32]
  wire [31:0] binaryOp_mul5762_io_Out_0_bits_data; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_io_LeftIO_ready; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_io_LeftIO_valid; // @[extracted_function_conv.scala 275:32]
  wire [31:0] binaryOp_mul5762_io_LeftIO_bits_data; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_io_RightIO_ready; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_mul5762_io_RightIO_valid; // @[extracted_function_conv.scala 275:32]
  wire [31:0] binaryOp_mul5762_io_RightIO_bits_data; // @[extracted_function_conv.scala 275:32]
  wire  binaryOp_add5863_clock; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_reset; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_enable_ready; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_enable_valid; // @[extracted_function_conv.scala 278:32]
  wire [4:0] binaryOp_add5863_io_enable_bits_taskID; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_enable_bits_control; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_Out_0_ready; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_Out_0_valid; // @[extracted_function_conv.scala 278:32]
  wire [4:0] binaryOp_add5863_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 278:32]
  wire [31:0] binaryOp_add5863_io_Out_0_bits_data; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_Out_1_ready; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_Out_1_valid; // @[extracted_function_conv.scala 278:32]
  wire [31:0] binaryOp_add5863_io_Out_1_bits_data; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_LeftIO_ready; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_LeftIO_valid; // @[extracted_function_conv.scala 278:32]
  wire [31:0] binaryOp_add5863_io_LeftIO_bits_data; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_RightIO_ready; // @[extracted_function_conv.scala 278:32]
  wire  binaryOp_add5863_io_RightIO_valid; // @[extracted_function_conv.scala 278:32]
  wire [31:0] binaryOp_add5863_io_RightIO_bits_data; // @[extracted_function_conv.scala 278:32]
  wire  st_64_clock; // @[extracted_function_conv.scala 281:21]
  wire  st_64_reset; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_enable_ready; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_enable_valid; // @[extracted_function_conv.scala 281:21]
  wire [4:0] st_64_io_enable_bits_taskID; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_enable_bits_control; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_GepAddr_ready; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_GepAddr_valid; // @[extracted_function_conv.scala 281:21]
  wire [4:0] st_64_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 281:21]
  wire [31:0] st_64_io_GepAddr_bits_data; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_inData_ready; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_inData_valid; // @[extracted_function_conv.scala 281:21]
  wire [4:0] st_64_io_inData_bits_taskID; // @[extracted_function_conv.scala 281:21]
  wire [31:0] st_64_io_inData_bits_data; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_memReq_ready; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_memReq_valid; // @[extracted_function_conv.scala 281:21]
  wire [21:0] st_64_io_memReq_bits_address; // @[extracted_function_conv.scala 281:21]
  wire [31:0] st_64_io_memReq_bits_data; // @[extracted_function_conv.scala 281:21]
  wire [4:0] st_64_io_memReq_bits_taskID; // @[extracted_function_conv.scala 281:21]
  wire  st_64_io_memResp_valid; // @[extracted_function_conv.scala 281:21]
  wire  ld_65_clock; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_reset; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_enable_ready; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_enable_valid; // @[extracted_function_conv.scala 284:21]
  wire [4:0] ld_65_io_enable_bits_taskID; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_enable_bits_control; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_Out_0_ready; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_Out_0_valid; // @[extracted_function_conv.scala 284:21]
  wire [31:0] ld_65_io_Out_0_bits_data; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_GepAddr_ready; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_GepAddr_valid; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 284:21]
  wire [4:0] ld_65_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 284:21]
  wire [31:0] ld_65_io_GepAddr_bits_data; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_memReq_ready; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_memReq_valid; // @[extracted_function_conv.scala 284:21]
  wire [31:0] ld_65_io_memReq_bits_address; // @[extracted_function_conv.scala 284:21]
  wire [4:0] ld_65_io_memReq_bits_taskID; // @[extracted_function_conv.scala 284:21]
  wire  ld_65_io_memResp_valid; // @[extracted_function_conv.scala 284:21]
  wire [31:0] ld_65_io_memResp_data; // @[extracted_function_conv.scala 284:21]
  wire  binaryOp_add6566_clock; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_reset; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_io_enable_ready; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_io_enable_valid; // @[extracted_function_conv.scala 287:32]
  wire [4:0] binaryOp_add6566_io_enable_bits_taskID; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_io_enable_bits_control; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_io_Out_0_ready; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_io_Out_0_valid; // @[extracted_function_conv.scala 287:32]
  wire [31:0] binaryOp_add6566_io_Out_0_bits_data; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_io_LeftIO_ready; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_io_LeftIO_valid; // @[extracted_function_conv.scala 287:32]
  wire [31:0] binaryOp_add6566_io_LeftIO_bits_data; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_io_RightIO_ready; // @[extracted_function_conv.scala 287:32]
  wire  binaryOp_add6566_io_RightIO_valid; // @[extracted_function_conv.scala 287:32]
  wire  Gep_arrayidx6667_clock; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_reset; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_enable_ready; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_enable_valid; // @[extracted_function_conv.scala 290:32]
  wire [4:0] Gep_arrayidx6667_io_enable_bits_taskID; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_enable_bits_control; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_Out_0_ready; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_Out_0_valid; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 290:32]
  wire [4:0] Gep_arrayidx6667_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 290:32]
  wire [31:0] Gep_arrayidx6667_io_Out_0_bits_data; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_baseAddress_ready; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_baseAddress_valid; // @[extracted_function_conv.scala 290:32]
  wire [4:0] Gep_arrayidx6667_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 290:32]
  wire [31:0] Gep_arrayidx6667_io_baseAddress_bits_data; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_idx_0_ready; // @[extracted_function_conv.scala 290:32]
  wire  Gep_arrayidx6667_io_idx_0_valid; // @[extracted_function_conv.scala 290:32]
  wire [31:0] Gep_arrayidx6667_io_idx_0_bits_data; // @[extracted_function_conv.scala 290:32]
  wire  ld_68_clock; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_reset; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_enable_ready; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_enable_valid; // @[extracted_function_conv.scala 293:21]
  wire [4:0] ld_68_io_enable_bits_taskID; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_enable_bits_control; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_Out_0_ready; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_Out_0_valid; // @[extracted_function_conv.scala 293:21]
  wire [31:0] ld_68_io_Out_0_bits_data; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_GepAddr_ready; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_GepAddr_valid; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 293:21]
  wire [4:0] ld_68_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 293:21]
  wire [31:0] ld_68_io_GepAddr_bits_data; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_memReq_ready; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_memReq_valid; // @[extracted_function_conv.scala 293:21]
  wire [31:0] ld_68_io_memReq_bits_address; // @[extracted_function_conv.scala 293:21]
  wire [4:0] ld_68_io_memReq_bits_taskID; // @[extracted_function_conv.scala 293:21]
  wire  ld_68_io_memResp_valid; // @[extracted_function_conv.scala 293:21]
  wire [31:0] ld_68_io_memResp_data; // @[extracted_function_conv.scala 293:21]
  wire  sextconv6869_clock; // @[extracted_function_conv.scala 296:28]
  wire  sextconv6869_reset; // @[extracted_function_conv.scala 296:28]
  wire  sextconv6869_io_Input_ready; // @[extracted_function_conv.scala 296:28]
  wire  sextconv6869_io_Input_valid; // @[extracted_function_conv.scala 296:28]
  wire [31:0] sextconv6869_io_Input_bits_data; // @[extracted_function_conv.scala 296:28]
  wire  sextconv6869_io_enable_ready; // @[extracted_function_conv.scala 296:28]
  wire  sextconv6869_io_enable_valid; // @[extracted_function_conv.scala 296:28]
  wire [4:0] sextconv6869_io_enable_bits_taskID; // @[extracted_function_conv.scala 296:28]
  wire  sextconv6869_io_Out_0_ready; // @[extracted_function_conv.scala 296:28]
  wire  sextconv6869_io_Out_0_valid; // @[extracted_function_conv.scala 296:28]
  wire [31:0] sextconv6869_io_Out_0_bits_data; // @[extracted_function_conv.scala 296:28]
  wire  binaryOp_mul6970_clock; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_reset; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_io_enable_ready; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_io_enable_valid; // @[extracted_function_conv.scala 299:32]
  wire [4:0] binaryOp_mul6970_io_enable_bits_taskID; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_io_enable_bits_control; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_io_Out_0_ready; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_io_Out_0_valid; // @[extracted_function_conv.scala 299:32]
  wire [31:0] binaryOp_mul6970_io_Out_0_bits_data; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_io_LeftIO_ready; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_io_LeftIO_valid; // @[extracted_function_conv.scala 299:32]
  wire [31:0] binaryOp_mul6970_io_LeftIO_bits_data; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_io_RightIO_ready; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_mul6970_io_RightIO_valid; // @[extracted_function_conv.scala 299:32]
  wire [31:0] binaryOp_mul6970_io_RightIO_bits_data; // @[extracted_function_conv.scala 299:32]
  wire  binaryOp_add7071_clock; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_reset; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_enable_ready; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_enable_valid; // @[extracted_function_conv.scala 302:32]
  wire [4:0] binaryOp_add7071_io_enable_bits_taskID; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_enable_bits_control; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_Out_0_ready; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_Out_0_valid; // @[extracted_function_conv.scala 302:32]
  wire [4:0] binaryOp_add7071_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 302:32]
  wire [31:0] binaryOp_add7071_io_Out_0_bits_data; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_Out_1_ready; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_Out_1_valid; // @[extracted_function_conv.scala 302:32]
  wire [31:0] binaryOp_add7071_io_Out_1_bits_data; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_LeftIO_ready; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_LeftIO_valid; // @[extracted_function_conv.scala 302:32]
  wire [31:0] binaryOp_add7071_io_LeftIO_bits_data; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_RightIO_ready; // @[extracted_function_conv.scala 302:32]
  wire  binaryOp_add7071_io_RightIO_valid; // @[extracted_function_conv.scala 302:32]
  wire [31:0] binaryOp_add7071_io_RightIO_bits_data; // @[extracted_function_conv.scala 302:32]
  wire  st_72_clock; // @[extracted_function_conv.scala 305:21]
  wire  st_72_reset; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_enable_ready; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_enable_valid; // @[extracted_function_conv.scala 305:21]
  wire [4:0] st_72_io_enable_bits_taskID; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_enable_bits_control; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_GepAddr_ready; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_GepAddr_valid; // @[extracted_function_conv.scala 305:21]
  wire [4:0] st_72_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 305:21]
  wire [31:0] st_72_io_GepAddr_bits_data; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_inData_ready; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_inData_valid; // @[extracted_function_conv.scala 305:21]
  wire [4:0] st_72_io_inData_bits_taskID; // @[extracted_function_conv.scala 305:21]
  wire [31:0] st_72_io_inData_bits_data; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_memReq_ready; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_memReq_valid; // @[extracted_function_conv.scala 305:21]
  wire [21:0] st_72_io_memReq_bits_address; // @[extracted_function_conv.scala 305:21]
  wire [31:0] st_72_io_memReq_bits_data; // @[extracted_function_conv.scala 305:21]
  wire [4:0] st_72_io_memReq_bits_taskID; // @[extracted_function_conv.scala 305:21]
  wire  st_72_io_memResp_valid; // @[extracted_function_conv.scala 305:21]
  wire  ld_73_clock; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_reset; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_enable_ready; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_enable_valid; // @[extracted_function_conv.scala 308:21]
  wire [4:0] ld_73_io_enable_bits_taskID; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_enable_bits_control; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_Out_0_ready; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_Out_0_valid; // @[extracted_function_conv.scala 308:21]
  wire [31:0] ld_73_io_Out_0_bits_data; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_GepAddr_ready; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_GepAddr_valid; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 308:21]
  wire [4:0] ld_73_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 308:21]
  wire [31:0] ld_73_io_GepAddr_bits_data; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_memReq_ready; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_memReq_valid; // @[extracted_function_conv.scala 308:21]
  wire [31:0] ld_73_io_memReq_bits_address; // @[extracted_function_conv.scala 308:21]
  wire [4:0] ld_73_io_memReq_bits_taskID; // @[extracted_function_conv.scala 308:21]
  wire  ld_73_io_memResp_valid; // @[extracted_function_conv.scala 308:21]
  wire [31:0] ld_73_io_memResp_data; // @[extracted_function_conv.scala 308:21]
  wire  binaryOp_add7774_clock; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_reset; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_io_enable_ready; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_io_enable_valid; // @[extracted_function_conv.scala 311:32]
  wire [4:0] binaryOp_add7774_io_enable_bits_taskID; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_io_enable_bits_control; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_io_Out_0_ready; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_io_Out_0_valid; // @[extracted_function_conv.scala 311:32]
  wire [31:0] binaryOp_add7774_io_Out_0_bits_data; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_io_LeftIO_ready; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_io_LeftIO_valid; // @[extracted_function_conv.scala 311:32]
  wire [31:0] binaryOp_add7774_io_LeftIO_bits_data; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_io_RightIO_ready; // @[extracted_function_conv.scala 311:32]
  wire  binaryOp_add7774_io_RightIO_valid; // @[extracted_function_conv.scala 311:32]
  wire  Gep_arrayidx7875_clock; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_reset; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_enable_ready; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_enable_valid; // @[extracted_function_conv.scala 314:32]
  wire [4:0] Gep_arrayidx7875_io_enable_bits_taskID; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_enable_bits_control; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_Out_0_ready; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_Out_0_valid; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 314:32]
  wire [4:0] Gep_arrayidx7875_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 314:32]
  wire [31:0] Gep_arrayidx7875_io_Out_0_bits_data; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_baseAddress_ready; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_baseAddress_valid; // @[extracted_function_conv.scala 314:32]
  wire [4:0] Gep_arrayidx7875_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 314:32]
  wire [31:0] Gep_arrayidx7875_io_baseAddress_bits_data; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_idx_0_ready; // @[extracted_function_conv.scala 314:32]
  wire  Gep_arrayidx7875_io_idx_0_valid; // @[extracted_function_conv.scala 314:32]
  wire [31:0] Gep_arrayidx7875_io_idx_0_bits_data; // @[extracted_function_conv.scala 314:32]
  wire  ld_76_clock; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_reset; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_enable_ready; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_enable_valid; // @[extracted_function_conv.scala 317:21]
  wire [4:0] ld_76_io_enable_bits_taskID; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_enable_bits_control; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_Out_0_ready; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_Out_0_valid; // @[extracted_function_conv.scala 317:21]
  wire [31:0] ld_76_io_Out_0_bits_data; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_GepAddr_ready; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_GepAddr_valid; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 317:21]
  wire [4:0] ld_76_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 317:21]
  wire [31:0] ld_76_io_GepAddr_bits_data; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_memReq_ready; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_memReq_valid; // @[extracted_function_conv.scala 317:21]
  wire [31:0] ld_76_io_memReq_bits_address; // @[extracted_function_conv.scala 317:21]
  wire [4:0] ld_76_io_memReq_bits_taskID; // @[extracted_function_conv.scala 317:21]
  wire  ld_76_io_memResp_valid; // @[extracted_function_conv.scala 317:21]
  wire [31:0] ld_76_io_memResp_data; // @[extracted_function_conv.scala 317:21]
  wire  sextconv8077_clock; // @[extracted_function_conv.scala 320:28]
  wire  sextconv8077_reset; // @[extracted_function_conv.scala 320:28]
  wire  sextconv8077_io_Input_ready; // @[extracted_function_conv.scala 320:28]
  wire  sextconv8077_io_Input_valid; // @[extracted_function_conv.scala 320:28]
  wire [31:0] sextconv8077_io_Input_bits_data; // @[extracted_function_conv.scala 320:28]
  wire  sextconv8077_io_enable_ready; // @[extracted_function_conv.scala 320:28]
  wire  sextconv8077_io_enable_valid; // @[extracted_function_conv.scala 320:28]
  wire [4:0] sextconv8077_io_enable_bits_taskID; // @[extracted_function_conv.scala 320:28]
  wire  sextconv8077_io_Out_0_ready; // @[extracted_function_conv.scala 320:28]
  wire  sextconv8077_io_Out_0_valid; // @[extracted_function_conv.scala 320:28]
  wire [31:0] sextconv8077_io_Out_0_bits_data; // @[extracted_function_conv.scala 320:28]
  wire  binaryOp_mul8178_clock; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_reset; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_io_enable_ready; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_io_enable_valid; // @[extracted_function_conv.scala 323:32]
  wire [4:0] binaryOp_mul8178_io_enable_bits_taskID; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_io_enable_bits_control; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_io_Out_0_ready; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_io_Out_0_valid; // @[extracted_function_conv.scala 323:32]
  wire [31:0] binaryOp_mul8178_io_Out_0_bits_data; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_io_LeftIO_ready; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_io_LeftIO_valid; // @[extracted_function_conv.scala 323:32]
  wire [31:0] binaryOp_mul8178_io_LeftIO_bits_data; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_io_RightIO_ready; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_mul8178_io_RightIO_valid; // @[extracted_function_conv.scala 323:32]
  wire [31:0] binaryOp_mul8178_io_RightIO_bits_data; // @[extracted_function_conv.scala 323:32]
  wire  binaryOp_add8279_clock; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_reset; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_enable_ready; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_enable_valid; // @[extracted_function_conv.scala 326:32]
  wire [4:0] binaryOp_add8279_io_enable_bits_taskID; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_enable_bits_control; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_Out_0_ready; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_Out_0_valid; // @[extracted_function_conv.scala 326:32]
  wire [4:0] binaryOp_add8279_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 326:32]
  wire [31:0] binaryOp_add8279_io_Out_0_bits_data; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_Out_1_ready; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_Out_1_valid; // @[extracted_function_conv.scala 326:32]
  wire [31:0] binaryOp_add8279_io_Out_1_bits_data; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_LeftIO_ready; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_LeftIO_valid; // @[extracted_function_conv.scala 326:32]
  wire [31:0] binaryOp_add8279_io_LeftIO_bits_data; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_RightIO_ready; // @[extracted_function_conv.scala 326:32]
  wire  binaryOp_add8279_io_RightIO_valid; // @[extracted_function_conv.scala 326:32]
  wire [31:0] binaryOp_add8279_io_RightIO_bits_data; // @[extracted_function_conv.scala 326:32]
  wire  st_80_clock; // @[extracted_function_conv.scala 329:21]
  wire  st_80_reset; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_enable_ready; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_enable_valid; // @[extracted_function_conv.scala 329:21]
  wire [4:0] st_80_io_enable_bits_taskID; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_enable_bits_control; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_GepAddr_ready; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_GepAddr_valid; // @[extracted_function_conv.scala 329:21]
  wire [4:0] st_80_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 329:21]
  wire [31:0] st_80_io_GepAddr_bits_data; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_inData_ready; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_inData_valid; // @[extracted_function_conv.scala 329:21]
  wire [4:0] st_80_io_inData_bits_taskID; // @[extracted_function_conv.scala 329:21]
  wire [31:0] st_80_io_inData_bits_data; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_memReq_ready; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_memReq_valid; // @[extracted_function_conv.scala 329:21]
  wire [21:0] st_80_io_memReq_bits_address; // @[extracted_function_conv.scala 329:21]
  wire [31:0] st_80_io_memReq_bits_data; // @[extracted_function_conv.scala 329:21]
  wire [4:0] st_80_io_memReq_bits_taskID; // @[extracted_function_conv.scala 329:21]
  wire  st_80_io_memResp_valid; // @[extracted_function_conv.scala 329:21]
  wire  ld_81_clock; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_reset; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_enable_ready; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_enable_valid; // @[extracted_function_conv.scala 332:21]
  wire [4:0] ld_81_io_enable_bits_taskID; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_enable_bits_control; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_Out_0_ready; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_Out_0_valid; // @[extracted_function_conv.scala 332:21]
  wire [31:0] ld_81_io_Out_0_bits_data; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_GepAddr_ready; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_GepAddr_valid; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 332:21]
  wire [4:0] ld_81_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 332:21]
  wire [31:0] ld_81_io_GepAddr_bits_data; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_memReq_ready; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_memReq_valid; // @[extracted_function_conv.scala 332:21]
  wire [31:0] ld_81_io_memReq_bits_address; // @[extracted_function_conv.scala 332:21]
  wire [4:0] ld_81_io_memReq_bits_taskID; // @[extracted_function_conv.scala 332:21]
  wire  ld_81_io_memResp_valid; // @[extracted_function_conv.scala 332:21]
  wire [31:0] ld_81_io_memResp_data; // @[extracted_function_conv.scala 332:21]
  wire  binaryOp_add8882_clock; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_reset; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_enable_ready; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_enable_valid; // @[extracted_function_conv.scala 335:32]
  wire [4:0] binaryOp_add8882_io_enable_bits_taskID; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_enable_bits_control; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_Out_0_ready; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_Out_0_valid; // @[extracted_function_conv.scala 335:32]
  wire [31:0] binaryOp_add8882_io_Out_0_bits_data; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_Out_1_ready; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_Out_1_valid; // @[extracted_function_conv.scala 335:32]
  wire [31:0] binaryOp_add8882_io_Out_1_bits_data; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_Out_2_ready; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_Out_2_valid; // @[extracted_function_conv.scala 335:32]
  wire [31:0] binaryOp_add8882_io_Out_2_bits_data; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_LeftIO_ready; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_LeftIO_valid; // @[extracted_function_conv.scala 335:32]
  wire [31:0] binaryOp_add8882_io_LeftIO_bits_data; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_RightIO_ready; // @[extracted_function_conv.scala 335:32]
  wire  binaryOp_add8882_io_RightIO_valid; // @[extracted_function_conv.scala 335:32]
  wire [31:0] binaryOp_add8882_io_RightIO_bits_data; // @[extracted_function_conv.scala 335:32]
  wire  Gep_arrayidx8983_clock; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_reset; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_enable_ready; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_enable_valid; // @[extracted_function_conv.scala 338:32]
  wire [4:0] Gep_arrayidx8983_io_enable_bits_taskID; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_enable_bits_control; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_Out_0_ready; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_Out_0_valid; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 338:32]
  wire [4:0] Gep_arrayidx8983_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 338:32]
  wire [31:0] Gep_arrayidx8983_io_Out_0_bits_data; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_baseAddress_ready; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_baseAddress_valid; // @[extracted_function_conv.scala 338:32]
  wire [4:0] Gep_arrayidx8983_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 338:32]
  wire [31:0] Gep_arrayidx8983_io_baseAddress_bits_data; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_idx_0_ready; // @[extracted_function_conv.scala 338:32]
  wire  Gep_arrayidx8983_io_idx_0_valid; // @[extracted_function_conv.scala 338:32]
  wire [31:0] Gep_arrayidx8983_io_idx_0_bits_data; // @[extracted_function_conv.scala 338:32]
  wire  ld_84_clock; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_reset; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_enable_ready; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_enable_valid; // @[extracted_function_conv.scala 341:21]
  wire [4:0] ld_84_io_enable_bits_taskID; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_enable_bits_control; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_Out_0_ready; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_Out_0_valid; // @[extracted_function_conv.scala 341:21]
  wire [31:0] ld_84_io_Out_0_bits_data; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_GepAddr_ready; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_GepAddr_valid; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 341:21]
  wire [4:0] ld_84_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 341:21]
  wire [31:0] ld_84_io_GepAddr_bits_data; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_memReq_ready; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_memReq_valid; // @[extracted_function_conv.scala 341:21]
  wire [31:0] ld_84_io_memReq_bits_address; // @[extracted_function_conv.scala 341:21]
  wire [4:0] ld_84_io_memReq_bits_taskID; // @[extracted_function_conv.scala 341:21]
  wire  ld_84_io_memResp_valid; // @[extracted_function_conv.scala 341:21]
  wire [31:0] ld_84_io_memResp_data; // @[extracted_function_conv.scala 341:21]
  wire  sextconv9185_clock; // @[extracted_function_conv.scala 344:28]
  wire  sextconv9185_reset; // @[extracted_function_conv.scala 344:28]
  wire  sextconv9185_io_Input_ready; // @[extracted_function_conv.scala 344:28]
  wire  sextconv9185_io_Input_valid; // @[extracted_function_conv.scala 344:28]
  wire [31:0] sextconv9185_io_Input_bits_data; // @[extracted_function_conv.scala 344:28]
  wire  sextconv9185_io_enable_ready; // @[extracted_function_conv.scala 344:28]
  wire  sextconv9185_io_enable_valid; // @[extracted_function_conv.scala 344:28]
  wire [4:0] sextconv9185_io_enable_bits_taskID; // @[extracted_function_conv.scala 344:28]
  wire  sextconv9185_io_Out_0_ready; // @[extracted_function_conv.scala 344:28]
  wire  sextconv9185_io_Out_0_valid; // @[extracted_function_conv.scala 344:28]
  wire [31:0] sextconv9185_io_Out_0_bits_data; // @[extracted_function_conv.scala 344:28]
  wire  binaryOp_mul9286_clock; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_reset; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_io_enable_ready; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_io_enable_valid; // @[extracted_function_conv.scala 347:32]
  wire [4:0] binaryOp_mul9286_io_enable_bits_taskID; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_io_enable_bits_control; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_io_Out_0_ready; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_io_Out_0_valid; // @[extracted_function_conv.scala 347:32]
  wire [31:0] binaryOp_mul9286_io_Out_0_bits_data; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_io_LeftIO_ready; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_io_LeftIO_valid; // @[extracted_function_conv.scala 347:32]
  wire [31:0] binaryOp_mul9286_io_LeftIO_bits_data; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_io_RightIO_ready; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_mul9286_io_RightIO_valid; // @[extracted_function_conv.scala 347:32]
  wire [31:0] binaryOp_mul9286_io_RightIO_bits_data; // @[extracted_function_conv.scala 347:32]
  wire  binaryOp_add9387_clock; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_reset; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_enable_ready; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_enable_valid; // @[extracted_function_conv.scala 350:32]
  wire [4:0] binaryOp_add9387_io_enable_bits_taskID; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_enable_bits_control; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_Out_0_ready; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_Out_0_valid; // @[extracted_function_conv.scala 350:32]
  wire [4:0] binaryOp_add9387_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 350:32]
  wire [31:0] binaryOp_add9387_io_Out_0_bits_data; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_Out_1_ready; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_Out_1_valid; // @[extracted_function_conv.scala 350:32]
  wire [31:0] binaryOp_add9387_io_Out_1_bits_data; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_LeftIO_ready; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_LeftIO_valid; // @[extracted_function_conv.scala 350:32]
  wire [31:0] binaryOp_add9387_io_LeftIO_bits_data; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_RightIO_ready; // @[extracted_function_conv.scala 350:32]
  wire  binaryOp_add9387_io_RightIO_valid; // @[extracted_function_conv.scala 350:32]
  wire [31:0] binaryOp_add9387_io_RightIO_bits_data; // @[extracted_function_conv.scala 350:32]
  wire  st_88_clock; // @[extracted_function_conv.scala 353:21]
  wire  st_88_reset; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_enable_ready; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_enable_valid; // @[extracted_function_conv.scala 353:21]
  wire [4:0] st_88_io_enable_bits_taskID; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_enable_bits_control; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_GepAddr_ready; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_GepAddr_valid; // @[extracted_function_conv.scala 353:21]
  wire [4:0] st_88_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 353:21]
  wire [31:0] st_88_io_GepAddr_bits_data; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_inData_ready; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_inData_valid; // @[extracted_function_conv.scala 353:21]
  wire [4:0] st_88_io_inData_bits_taskID; // @[extracted_function_conv.scala 353:21]
  wire [31:0] st_88_io_inData_bits_data; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_memReq_ready; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_memReq_valid; // @[extracted_function_conv.scala 353:21]
  wire [21:0] st_88_io_memReq_bits_address; // @[extracted_function_conv.scala 353:21]
  wire [31:0] st_88_io_memReq_bits_data; // @[extracted_function_conv.scala 353:21]
  wire [4:0] st_88_io_memReq_bits_taskID; // @[extracted_function_conv.scala 353:21]
  wire  st_88_io_memResp_valid; // @[extracted_function_conv.scala 353:21]
  wire  ld_89_clock; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_reset; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_enable_ready; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_enable_valid; // @[extracted_function_conv.scala 356:21]
  wire [4:0] ld_89_io_enable_bits_taskID; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_enable_bits_control; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_Out_0_ready; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_Out_0_valid; // @[extracted_function_conv.scala 356:21]
  wire [31:0] ld_89_io_Out_0_bits_data; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_GepAddr_ready; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_GepAddr_valid; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 356:21]
  wire [4:0] ld_89_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 356:21]
  wire [31:0] ld_89_io_GepAddr_bits_data; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_memReq_ready; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_memReq_valid; // @[extracted_function_conv.scala 356:21]
  wire [31:0] ld_89_io_memReq_bits_address; // @[extracted_function_conv.scala 356:21]
  wire [4:0] ld_89_io_memReq_bits_taskID; // @[extracted_function_conv.scala 356:21]
  wire  ld_89_io_memResp_valid; // @[extracted_function_conv.scala 356:21]
  wire [31:0] ld_89_io_memResp_data; // @[extracted_function_conv.scala 356:21]
  wire  binaryOp_add10090_clock; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_reset; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_io_enable_ready; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_io_enable_valid; // @[extracted_function_conv.scala 359:33]
  wire [4:0] binaryOp_add10090_io_enable_bits_taskID; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_io_enable_bits_control; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_io_Out_0_ready; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_io_Out_0_valid; // @[extracted_function_conv.scala 359:33]
  wire [31:0] binaryOp_add10090_io_Out_0_bits_data; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_io_LeftIO_ready; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_io_LeftIO_valid; // @[extracted_function_conv.scala 359:33]
  wire [31:0] binaryOp_add10090_io_LeftIO_bits_data; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_io_RightIO_ready; // @[extracted_function_conv.scala 359:33]
  wire  binaryOp_add10090_io_RightIO_valid; // @[extracted_function_conv.scala 359:33]
  wire  Gep_arrayidx10191_clock; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_reset; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_enable_ready; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_enable_valid; // @[extracted_function_conv.scala 362:33]
  wire [4:0] Gep_arrayidx10191_io_enable_bits_taskID; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_enable_bits_control; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_Out_0_ready; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_Out_0_valid; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 362:33]
  wire [4:0] Gep_arrayidx10191_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 362:33]
  wire [31:0] Gep_arrayidx10191_io_Out_0_bits_data; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_baseAddress_ready; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_baseAddress_valid; // @[extracted_function_conv.scala 362:33]
  wire [4:0] Gep_arrayidx10191_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 362:33]
  wire [31:0] Gep_arrayidx10191_io_baseAddress_bits_data; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_idx_0_ready; // @[extracted_function_conv.scala 362:33]
  wire  Gep_arrayidx10191_io_idx_0_valid; // @[extracted_function_conv.scala 362:33]
  wire [31:0] Gep_arrayidx10191_io_idx_0_bits_data; // @[extracted_function_conv.scala 362:33]
  wire  ld_92_clock; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_reset; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_enable_ready; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_enable_valid; // @[extracted_function_conv.scala 365:21]
  wire [4:0] ld_92_io_enable_bits_taskID; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_enable_bits_control; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_Out_0_ready; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_Out_0_valid; // @[extracted_function_conv.scala 365:21]
  wire [31:0] ld_92_io_Out_0_bits_data; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_GepAddr_ready; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_GepAddr_valid; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 365:21]
  wire [4:0] ld_92_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 365:21]
  wire [31:0] ld_92_io_GepAddr_bits_data; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_memReq_ready; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_memReq_valid; // @[extracted_function_conv.scala 365:21]
  wire [31:0] ld_92_io_memReq_bits_address; // @[extracted_function_conv.scala 365:21]
  wire [4:0] ld_92_io_memReq_bits_taskID; // @[extracted_function_conv.scala 365:21]
  wire  ld_92_io_memResp_valid; // @[extracted_function_conv.scala 365:21]
  wire [31:0] ld_92_io_memResp_data; // @[extracted_function_conv.scala 365:21]
  wire  sextconv10393_clock; // @[extracted_function_conv.scala 368:29]
  wire  sextconv10393_reset; // @[extracted_function_conv.scala 368:29]
  wire  sextconv10393_io_Input_ready; // @[extracted_function_conv.scala 368:29]
  wire  sextconv10393_io_Input_valid; // @[extracted_function_conv.scala 368:29]
  wire [31:0] sextconv10393_io_Input_bits_data; // @[extracted_function_conv.scala 368:29]
  wire  sextconv10393_io_enable_ready; // @[extracted_function_conv.scala 368:29]
  wire  sextconv10393_io_enable_valid; // @[extracted_function_conv.scala 368:29]
  wire [4:0] sextconv10393_io_enable_bits_taskID; // @[extracted_function_conv.scala 368:29]
  wire  sextconv10393_io_Out_0_ready; // @[extracted_function_conv.scala 368:29]
  wire  sextconv10393_io_Out_0_valid; // @[extracted_function_conv.scala 368:29]
  wire [31:0] sextconv10393_io_Out_0_bits_data; // @[extracted_function_conv.scala 368:29]
  wire  binaryOp_mul10494_clock; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_reset; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_io_enable_ready; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_io_enable_valid; // @[extracted_function_conv.scala 371:33]
  wire [4:0] binaryOp_mul10494_io_enable_bits_taskID; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_io_enable_bits_control; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_io_Out_0_ready; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_io_Out_0_valid; // @[extracted_function_conv.scala 371:33]
  wire [31:0] binaryOp_mul10494_io_Out_0_bits_data; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_io_LeftIO_ready; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_io_LeftIO_valid; // @[extracted_function_conv.scala 371:33]
  wire [31:0] binaryOp_mul10494_io_LeftIO_bits_data; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_io_RightIO_ready; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_mul10494_io_RightIO_valid; // @[extracted_function_conv.scala 371:33]
  wire [31:0] binaryOp_mul10494_io_RightIO_bits_data; // @[extracted_function_conv.scala 371:33]
  wire  binaryOp_add10595_clock; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_reset; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_enable_ready; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_enable_valid; // @[extracted_function_conv.scala 374:33]
  wire [4:0] binaryOp_add10595_io_enable_bits_taskID; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_enable_bits_control; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_Out_0_ready; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_Out_0_valid; // @[extracted_function_conv.scala 374:33]
  wire [4:0] binaryOp_add10595_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 374:33]
  wire [31:0] binaryOp_add10595_io_Out_0_bits_data; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_Out_1_ready; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_Out_1_valid; // @[extracted_function_conv.scala 374:33]
  wire [31:0] binaryOp_add10595_io_Out_1_bits_data; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_LeftIO_ready; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_LeftIO_valid; // @[extracted_function_conv.scala 374:33]
  wire [31:0] binaryOp_add10595_io_LeftIO_bits_data; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_RightIO_ready; // @[extracted_function_conv.scala 374:33]
  wire  binaryOp_add10595_io_RightIO_valid; // @[extracted_function_conv.scala 374:33]
  wire [31:0] binaryOp_add10595_io_RightIO_bits_data; // @[extracted_function_conv.scala 374:33]
  wire  st_96_clock; // @[extracted_function_conv.scala 377:21]
  wire  st_96_reset; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_enable_ready; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_enable_valid; // @[extracted_function_conv.scala 377:21]
  wire [4:0] st_96_io_enable_bits_taskID; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_enable_bits_control; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_GepAddr_ready; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_GepAddr_valid; // @[extracted_function_conv.scala 377:21]
  wire [4:0] st_96_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 377:21]
  wire [31:0] st_96_io_GepAddr_bits_data; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_inData_ready; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_inData_valid; // @[extracted_function_conv.scala 377:21]
  wire [4:0] st_96_io_inData_bits_taskID; // @[extracted_function_conv.scala 377:21]
  wire [31:0] st_96_io_inData_bits_data; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_memReq_ready; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_memReq_valid; // @[extracted_function_conv.scala 377:21]
  wire [21:0] st_96_io_memReq_bits_address; // @[extracted_function_conv.scala 377:21]
  wire [31:0] st_96_io_memReq_bits_data; // @[extracted_function_conv.scala 377:21]
  wire [4:0] st_96_io_memReq_bits_taskID; // @[extracted_function_conv.scala 377:21]
  wire  st_96_io_memResp_valid; // @[extracted_function_conv.scala 377:21]
  wire  ld_97_clock; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_reset; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_enable_ready; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_enable_valid; // @[extracted_function_conv.scala 380:21]
  wire [4:0] ld_97_io_enable_bits_taskID; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_enable_bits_control; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_Out_0_ready; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_Out_0_valid; // @[extracted_function_conv.scala 380:21]
  wire [31:0] ld_97_io_Out_0_bits_data; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_GepAddr_ready; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_GepAddr_valid; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 380:21]
  wire [4:0] ld_97_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 380:21]
  wire [31:0] ld_97_io_GepAddr_bits_data; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_memReq_ready; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_memReq_valid; // @[extracted_function_conv.scala 380:21]
  wire [31:0] ld_97_io_memReq_bits_address; // @[extracted_function_conv.scala 380:21]
  wire [4:0] ld_97_io_memReq_bits_taskID; // @[extracted_function_conv.scala 380:21]
  wire  ld_97_io_memResp_valid; // @[extracted_function_conv.scala 380:21]
  wire [31:0] ld_97_io_memResp_data; // @[extracted_function_conv.scala 380:21]
  wire  binaryOp_add11298_clock; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_reset; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_io_enable_ready; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_io_enable_valid; // @[extracted_function_conv.scala 383:33]
  wire [4:0] binaryOp_add11298_io_enable_bits_taskID; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_io_enable_bits_control; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_io_Out_0_ready; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_io_Out_0_valid; // @[extracted_function_conv.scala 383:33]
  wire [31:0] binaryOp_add11298_io_Out_0_bits_data; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_io_LeftIO_ready; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_io_LeftIO_valid; // @[extracted_function_conv.scala 383:33]
  wire [31:0] binaryOp_add11298_io_LeftIO_bits_data; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_io_RightIO_ready; // @[extracted_function_conv.scala 383:33]
  wire  binaryOp_add11298_io_RightIO_valid; // @[extracted_function_conv.scala 383:33]
  wire  Gep_arrayidx11399_clock; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_reset; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_enable_ready; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_enable_valid; // @[extracted_function_conv.scala 386:33]
  wire [4:0] Gep_arrayidx11399_io_enable_bits_taskID; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_enable_bits_control; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_Out_0_ready; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_Out_0_valid; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 386:33]
  wire [4:0] Gep_arrayidx11399_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 386:33]
  wire [31:0] Gep_arrayidx11399_io_Out_0_bits_data; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_baseAddress_ready; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_baseAddress_valid; // @[extracted_function_conv.scala 386:33]
  wire [4:0] Gep_arrayidx11399_io_baseAddress_bits_taskID; // @[extracted_function_conv.scala 386:33]
  wire [31:0] Gep_arrayidx11399_io_baseAddress_bits_data; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_idx_0_ready; // @[extracted_function_conv.scala 386:33]
  wire  Gep_arrayidx11399_io_idx_0_valid; // @[extracted_function_conv.scala 386:33]
  wire [31:0] Gep_arrayidx11399_io_idx_0_bits_data; // @[extracted_function_conv.scala 386:33]
  wire  ld_100_clock; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_reset; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_enable_ready; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_enable_valid; // @[extracted_function_conv.scala 389:22]
  wire [4:0] ld_100_io_enable_bits_taskID; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_enable_bits_control; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_Out_0_ready; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_Out_0_valid; // @[extracted_function_conv.scala 389:22]
  wire [31:0] ld_100_io_Out_0_bits_data; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_GepAddr_ready; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_GepAddr_valid; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_GepAddr_bits_predicate; // @[extracted_function_conv.scala 389:22]
  wire [4:0] ld_100_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 389:22]
  wire [31:0] ld_100_io_GepAddr_bits_data; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_memReq_ready; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_memReq_valid; // @[extracted_function_conv.scala 389:22]
  wire [31:0] ld_100_io_memReq_bits_address; // @[extracted_function_conv.scala 389:22]
  wire [4:0] ld_100_io_memReq_bits_taskID; // @[extracted_function_conv.scala 389:22]
  wire  ld_100_io_memResp_valid; // @[extracted_function_conv.scala 389:22]
  wire [31:0] ld_100_io_memResp_data; // @[extracted_function_conv.scala 389:22]
  wire  sextconv115101_clock; // @[extracted_function_conv.scala 392:30]
  wire  sextconv115101_reset; // @[extracted_function_conv.scala 392:30]
  wire  sextconv115101_io_Input_ready; // @[extracted_function_conv.scala 392:30]
  wire  sextconv115101_io_Input_valid; // @[extracted_function_conv.scala 392:30]
  wire [31:0] sextconv115101_io_Input_bits_data; // @[extracted_function_conv.scala 392:30]
  wire  sextconv115101_io_enable_ready; // @[extracted_function_conv.scala 392:30]
  wire  sextconv115101_io_enable_valid; // @[extracted_function_conv.scala 392:30]
  wire [4:0] sextconv115101_io_enable_bits_taskID; // @[extracted_function_conv.scala 392:30]
  wire  sextconv115101_io_Out_0_ready; // @[extracted_function_conv.scala 392:30]
  wire  sextconv115101_io_Out_0_valid; // @[extracted_function_conv.scala 392:30]
  wire [31:0] sextconv115101_io_Out_0_bits_data; // @[extracted_function_conv.scala 392:30]
  wire  binaryOp_mul116102_clock; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_reset; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_io_enable_ready; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_io_enable_valid; // @[extracted_function_conv.scala 395:34]
  wire [4:0] binaryOp_mul116102_io_enable_bits_taskID; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_io_enable_bits_control; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_io_Out_0_ready; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_io_Out_0_valid; // @[extracted_function_conv.scala 395:34]
  wire [31:0] binaryOp_mul116102_io_Out_0_bits_data; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_io_LeftIO_ready; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_io_LeftIO_valid; // @[extracted_function_conv.scala 395:34]
  wire [31:0] binaryOp_mul116102_io_LeftIO_bits_data; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_io_RightIO_ready; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_mul116102_io_RightIO_valid; // @[extracted_function_conv.scala 395:34]
  wire [31:0] binaryOp_mul116102_io_RightIO_bits_data; // @[extracted_function_conv.scala 395:34]
  wire  binaryOp_add117103_clock; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_reset; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_io_enable_ready; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_io_enable_valid; // @[extracted_function_conv.scala 398:34]
  wire [4:0] binaryOp_add117103_io_enable_bits_taskID; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_io_enable_bits_control; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_io_Out_0_ready; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_io_Out_0_valid; // @[extracted_function_conv.scala 398:34]
  wire [4:0] binaryOp_add117103_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 398:34]
  wire [31:0] binaryOp_add117103_io_Out_0_bits_data; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_io_LeftIO_ready; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_io_LeftIO_valid; // @[extracted_function_conv.scala 398:34]
  wire [31:0] binaryOp_add117103_io_LeftIO_bits_data; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_io_RightIO_ready; // @[extracted_function_conv.scala 398:34]
  wire  binaryOp_add117103_io_RightIO_valid; // @[extracted_function_conv.scala 398:34]
  wire [31:0] binaryOp_add117103_io_RightIO_bits_data; // @[extracted_function_conv.scala 398:34]
  wire  st_104_clock; // @[extracted_function_conv.scala 401:22]
  wire  st_104_reset; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_enable_ready; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_enable_valid; // @[extracted_function_conv.scala 401:22]
  wire [4:0] st_104_io_enable_bits_taskID; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_enable_bits_control; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_GepAddr_ready; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_GepAddr_valid; // @[extracted_function_conv.scala 401:22]
  wire [4:0] st_104_io_GepAddr_bits_taskID; // @[extracted_function_conv.scala 401:22]
  wire [31:0] st_104_io_GepAddr_bits_data; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_inData_ready; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_inData_valid; // @[extracted_function_conv.scala 401:22]
  wire [4:0] st_104_io_inData_bits_taskID; // @[extracted_function_conv.scala 401:22]
  wire [31:0] st_104_io_inData_bits_data; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_memReq_ready; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_memReq_valid; // @[extracted_function_conv.scala 401:22]
  wire [21:0] st_104_io_memReq_bits_address; // @[extracted_function_conv.scala 401:22]
  wire [31:0] st_104_io_memReq_bits_data; // @[extracted_function_conv.scala 401:22]
  wire [4:0] st_104_io_memReq_bits_taskID; // @[extracted_function_conv.scala 401:22]
  wire  st_104_io_memResp_valid; // @[extracted_function_conv.scala 401:22]
  wire  binaryOp_inc105_clock; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_reset; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_enable_ready; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_enable_valid; // @[extracted_function_conv.scala 404:31]
  wire [4:0] binaryOp_inc105_io_enable_bits_taskID; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_enable_bits_control; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_Out_0_ready; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_Out_0_valid; // @[extracted_function_conv.scala 404:31]
  wire [4:0] binaryOp_inc105_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 404:31]
  wire [31:0] binaryOp_inc105_io_Out_0_bits_data; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_Out_1_ready; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_Out_1_valid; // @[extracted_function_conv.scala 404:31]
  wire [31:0] binaryOp_inc105_io_Out_1_bits_data; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_LeftIO_ready; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_LeftIO_valid; // @[extracted_function_conv.scala 404:31]
  wire [31:0] binaryOp_inc105_io_LeftIO_bits_data; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_RightIO_ready; // @[extracted_function_conv.scala 404:31]
  wire  binaryOp_inc105_io_RightIO_valid; // @[extracted_function_conv.scala 404:31]
  wire  icmp_exitcond106_clock; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_reset; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_io_enable_ready; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_io_enable_valid; // @[extracted_function_conv.scala 407:32]
  wire [4:0] icmp_exitcond106_io_enable_bits_taskID; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_io_enable_bits_control; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_io_Out_0_ready; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_io_Out_0_valid; // @[extracted_function_conv.scala 407:32]
  wire [4:0] icmp_exitcond106_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 407:32]
  wire [31:0] icmp_exitcond106_io_Out_0_bits_data; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_io_LeftIO_ready; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_io_LeftIO_valid; // @[extracted_function_conv.scala 407:32]
  wire [31:0] icmp_exitcond106_io_LeftIO_bits_data; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_io_RightIO_ready; // @[extracted_function_conv.scala 407:32]
  wire  icmp_exitcond106_io_RightIO_valid; // @[extracted_function_conv.scala 407:32]
  wire  br_107_clock; // @[extracted_function_conv.scala 410:22]
  wire  br_107_reset; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_enable_ready; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_enable_valid; // @[extracted_function_conv.scala 410:22]
  wire [4:0] br_107_io_enable_bits_taskID; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_enable_bits_control; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_CmpIO_ready; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_CmpIO_valid; // @[extracted_function_conv.scala 410:22]
  wire [4:0] br_107_io_CmpIO_bits_taskID; // @[extracted_function_conv.scala 410:22]
  wire [31:0] br_107_io_CmpIO_bits_data; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_TrueOutput_0_ready; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_TrueOutput_0_valid; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_TrueOutput_0_bits_control; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_FalseOutput_0_ready; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_FalseOutput_0_valid; // @[extracted_function_conv.scala 410:22]
  wire [4:0] br_107_io_FalseOutput_0_bits_taskID; // @[extracted_function_conv.scala 410:22]
  wire  br_107_io_FalseOutput_0_bits_control; // @[extracted_function_conv.scala 410:22]
  wire  const0_clock; // @[extracted_function_conv.scala 419:22]
  wire  const0_reset; // @[extracted_function_conv.scala 419:22]
  wire  const0_io_enable_ready; // @[extracted_function_conv.scala 419:22]
  wire  const0_io_enable_valid; // @[extracted_function_conv.scala 419:22]
  wire [4:0] const0_io_enable_bits_taskID; // @[extracted_function_conv.scala 419:22]
  wire  const0_io_Out_ready; // @[extracted_function_conv.scala 419:22]
  wire  const0_io_Out_valid; // @[extracted_function_conv.scala 419:22]
  wire  const1_clock; // @[extracted_function_conv.scala 422:22]
  wire  const1_reset; // @[extracted_function_conv.scala 422:22]
  wire  const1_io_enable_ready; // @[extracted_function_conv.scala 422:22]
  wire  const1_io_enable_valid; // @[extracted_function_conv.scala 422:22]
  wire [4:0] const1_io_enable_bits_taskID; // @[extracted_function_conv.scala 422:22]
  wire  const1_io_Out_ready; // @[extracted_function_conv.scala 422:22]
  wire  const1_io_Out_valid; // @[extracted_function_conv.scala 422:22]
  wire  const2_clock; // @[extracted_function_conv.scala 425:22]
  wire  const2_reset; // @[extracted_function_conv.scala 425:22]
  wire  const2_io_enable_ready; // @[extracted_function_conv.scala 425:22]
  wire  const2_io_enable_valid; // @[extracted_function_conv.scala 425:22]
  wire [4:0] const2_io_enable_bits_taskID; // @[extracted_function_conv.scala 425:22]
  wire  const2_io_Out_ready; // @[extracted_function_conv.scala 425:22]
  wire  const2_io_Out_valid; // @[extracted_function_conv.scala 425:22]
  wire  const3_clock; // @[extracted_function_conv.scala 428:22]
  wire  const3_reset; // @[extracted_function_conv.scala 428:22]
  wire  const3_io_enable_ready; // @[extracted_function_conv.scala 428:22]
  wire  const3_io_enable_valid; // @[extracted_function_conv.scala 428:22]
  wire [4:0] const3_io_enable_bits_taskID; // @[extracted_function_conv.scala 428:22]
  wire  const3_io_Out_ready; // @[extracted_function_conv.scala 428:22]
  wire  const3_io_Out_valid; // @[extracted_function_conv.scala 428:22]
  wire  const4_clock; // @[extracted_function_conv.scala 431:22]
  wire  const4_reset; // @[extracted_function_conv.scala 431:22]
  wire  const4_io_enable_ready; // @[extracted_function_conv.scala 431:22]
  wire  const4_io_enable_valid; // @[extracted_function_conv.scala 431:22]
  wire [4:0] const4_io_enable_bits_taskID; // @[extracted_function_conv.scala 431:22]
  wire  const4_io_Out_ready; // @[extracted_function_conv.scala 431:22]
  wire  const4_io_Out_valid; // @[extracted_function_conv.scala 431:22]
  wire  const5_clock; // @[extracted_function_conv.scala 434:22]
  wire  const5_reset; // @[extracted_function_conv.scala 434:22]
  wire  const5_io_enable_ready; // @[extracted_function_conv.scala 434:22]
  wire  const5_io_enable_valid; // @[extracted_function_conv.scala 434:22]
  wire [4:0] const5_io_enable_bits_taskID; // @[extracted_function_conv.scala 434:22]
  wire  const5_io_Out_ready; // @[extracted_function_conv.scala 434:22]
  wire  const5_io_Out_valid; // @[extracted_function_conv.scala 434:22]
  wire  const6_clock; // @[extracted_function_conv.scala 437:22]
  wire  const6_reset; // @[extracted_function_conv.scala 437:22]
  wire  const6_io_enable_ready; // @[extracted_function_conv.scala 437:22]
  wire  const6_io_enable_valid; // @[extracted_function_conv.scala 437:22]
  wire [4:0] const6_io_enable_bits_taskID; // @[extracted_function_conv.scala 437:22]
  wire  const6_io_Out_ready; // @[extracted_function_conv.scala 437:22]
  wire  const6_io_Out_valid; // @[extracted_function_conv.scala 437:22]
  wire  const7_clock; // @[extracted_function_conv.scala 440:22]
  wire  const7_reset; // @[extracted_function_conv.scala 440:22]
  wire  const7_io_enable_ready; // @[extracted_function_conv.scala 440:22]
  wire  const7_io_enable_valid; // @[extracted_function_conv.scala 440:22]
  wire [4:0] const7_io_enable_bits_taskID; // @[extracted_function_conv.scala 440:22]
  wire  const7_io_Out_ready; // @[extracted_function_conv.scala 440:22]
  wire  const7_io_Out_valid; // @[extracted_function_conv.scala 440:22]
  wire  const8_clock; // @[extracted_function_conv.scala 443:22]
  wire  const8_reset; // @[extracted_function_conv.scala 443:22]
  wire  const8_io_enable_ready; // @[extracted_function_conv.scala 443:22]
  wire  const8_io_enable_valid; // @[extracted_function_conv.scala 443:22]
  wire [4:0] const8_io_enable_bits_taskID; // @[extracted_function_conv.scala 443:22]
  wire  const8_io_Out_ready; // @[extracted_function_conv.scala 443:22]
  wire  const8_io_Out_valid; // @[extracted_function_conv.scala 443:22]
  wire [4:0] const8_io_Out_bits_taskID; // @[extracted_function_conv.scala 443:22]
  wire  const9_clock; // @[extracted_function_conv.scala 446:22]
  wire  const9_reset; // @[extracted_function_conv.scala 446:22]
  wire  const9_io_enable_ready; // @[extracted_function_conv.scala 446:22]
  wire  const9_io_enable_valid; // @[extracted_function_conv.scala 446:22]
  wire [4:0] const9_io_enable_bits_taskID; // @[extracted_function_conv.scala 446:22]
  wire  const9_io_Out_ready; // @[extracted_function_conv.scala 446:22]
  wire  const9_io_Out_valid; // @[extracted_function_conv.scala 446:22]
  wire  const10_clock; // @[extracted_function_conv.scala 449:23]
  wire  const10_reset; // @[extracted_function_conv.scala 449:23]
  wire  const10_io_enable_ready; // @[extracted_function_conv.scala 449:23]
  wire  const10_io_enable_valid; // @[extracted_function_conv.scala 449:23]
  wire [4:0] const10_io_enable_bits_taskID; // @[extracted_function_conv.scala 449:23]
  wire  const10_io_Out_ready; // @[extracted_function_conv.scala 449:23]
  wire  const10_io_Out_valid; // @[extracted_function_conv.scala 449:23]
  wire  const11_clock; // @[extracted_function_conv.scala 452:23]
  wire  const11_reset; // @[extracted_function_conv.scala 452:23]
  wire  const11_io_enable_ready; // @[extracted_function_conv.scala 452:23]
  wire  const11_io_enable_valid; // @[extracted_function_conv.scala 452:23]
  wire [4:0] const11_io_enable_bits_taskID; // @[extracted_function_conv.scala 452:23]
  wire  const11_io_Out_ready; // @[extracted_function_conv.scala 452:23]
  wire  const11_io_Out_valid; // @[extracted_function_conv.scala 452:23]
  wire  const12_clock; // @[extracted_function_conv.scala 455:23]
  wire  const12_reset; // @[extracted_function_conv.scala 455:23]
  wire  const12_io_enable_ready; // @[extracted_function_conv.scala 455:23]
  wire  const12_io_enable_valid; // @[extracted_function_conv.scala 455:23]
  wire [4:0] const12_io_enable_bits_taskID; // @[extracted_function_conv.scala 455:23]
  wire  const12_io_Out_ready; // @[extracted_function_conv.scala 455:23]
  wire  const12_io_Out_valid; // @[extracted_function_conv.scala 455:23]
  wire  const13_clock; // @[extracted_function_conv.scala 458:23]
  wire  const13_reset; // @[extracted_function_conv.scala 458:23]
  wire  const13_io_enable_ready; // @[extracted_function_conv.scala 458:23]
  wire  const13_io_enable_valid; // @[extracted_function_conv.scala 458:23]
  wire [4:0] const13_io_enable_bits_taskID; // @[extracted_function_conv.scala 458:23]
  wire  const13_io_Out_ready; // @[extracted_function_conv.scala 458:23]
  wire  const13_io_Out_valid; // @[extracted_function_conv.scala 458:23]
  wire  const14_clock; // @[extracted_function_conv.scala 461:23]
  wire  const14_reset; // @[extracted_function_conv.scala 461:23]
  wire  const14_io_enable_ready; // @[extracted_function_conv.scala 461:23]
  wire  const14_io_enable_valid; // @[extracted_function_conv.scala 461:23]
  wire [4:0] const14_io_enable_bits_taskID; // @[extracted_function_conv.scala 461:23]
  wire  const14_io_Out_ready; // @[extracted_function_conv.scala 461:23]
  wire  const14_io_Out_valid; // @[extracted_function_conv.scala 461:23]
  wire  const15_clock; // @[extracted_function_conv.scala 464:23]
  wire  const15_reset; // @[extracted_function_conv.scala 464:23]
  wire  const15_io_enable_ready; // @[extracted_function_conv.scala 464:23]
  wire  const15_io_enable_valid; // @[extracted_function_conv.scala 464:23]
  wire [4:0] const15_io_enable_bits_taskID; // @[extracted_function_conv.scala 464:23]
  wire  const15_io_Out_ready; // @[extracted_function_conv.scala 464:23]
  wire  const15_io_Out_valid; // @[extracted_function_conv.scala 464:23]
  wire [4:0] const15_io_Out_bits_taskID; // @[extracted_function_conv.scala 464:23]
  wire  const16_clock; // @[extracted_function_conv.scala 467:23]
  wire  const16_reset; // @[extracted_function_conv.scala 467:23]
  wire  const16_io_enable_ready; // @[extracted_function_conv.scala 467:23]
  wire  const16_io_enable_valid; // @[extracted_function_conv.scala 467:23]
  wire [4:0] const16_io_enable_bits_taskID; // @[extracted_function_conv.scala 467:23]
  wire  const16_io_Out_ready; // @[extracted_function_conv.scala 467:23]
  wire  const16_io_Out_valid; // @[extracted_function_conv.scala 467:23]
  wire  const17_clock; // @[extracted_function_conv.scala 470:23]
  wire  const17_reset; // @[extracted_function_conv.scala 470:23]
  wire  const17_io_enable_ready; // @[extracted_function_conv.scala 470:23]
  wire  const17_io_enable_valid; // @[extracted_function_conv.scala 470:23]
  wire [4:0] const17_io_enable_bits_taskID; // @[extracted_function_conv.scala 470:23]
  wire  const17_io_Out_ready; // @[extracted_function_conv.scala 470:23]
  wire  const17_io_Out_valid; // @[extracted_function_conv.scala 470:23]
  wire  const18_clock; // @[extracted_function_conv.scala 473:23]
  wire  const18_reset; // @[extracted_function_conv.scala 473:23]
  wire  const18_io_enable_ready; // @[extracted_function_conv.scala 473:23]
  wire  const18_io_enable_valid; // @[extracted_function_conv.scala 473:23]
  wire [4:0] const18_io_enable_bits_taskID; // @[extracted_function_conv.scala 473:23]
  wire  const18_io_Out_ready; // @[extracted_function_conv.scala 473:23]
  wire  const18_io_Out_valid; // @[extracted_function_conv.scala 473:23]
  wire  const19_clock; // @[extracted_function_conv.scala 476:23]
  wire  const19_reset; // @[extracted_function_conv.scala 476:23]
  wire  const19_io_enable_ready; // @[extracted_function_conv.scala 476:23]
  wire  const19_io_enable_valid; // @[extracted_function_conv.scala 476:23]
  wire [4:0] const19_io_enable_bits_taskID; // @[extracted_function_conv.scala 476:23]
  wire  const19_io_Out_ready; // @[extracted_function_conv.scala 476:23]
  wire  const19_io_Out_valid; // @[extracted_function_conv.scala 476:23]
  wire  const20_clock; // @[extracted_function_conv.scala 479:23]
  wire  const20_reset; // @[extracted_function_conv.scala 479:23]
  wire  const20_io_enable_ready; // @[extracted_function_conv.scala 479:23]
  wire  const20_io_enable_valid; // @[extracted_function_conv.scala 479:23]
  wire [4:0] const20_io_enable_bits_taskID; // @[extracted_function_conv.scala 479:23]
  wire  const20_io_Out_ready; // @[extracted_function_conv.scala 479:23]
  wire  const20_io_Out_valid; // @[extracted_function_conv.scala 479:23]
  wire  const21_clock; // @[extracted_function_conv.scala 482:23]
  wire  const21_reset; // @[extracted_function_conv.scala 482:23]
  wire  const21_io_enable_ready; // @[extracted_function_conv.scala 482:23]
  wire  const21_io_enable_valid; // @[extracted_function_conv.scala 482:23]
  wire [4:0] const21_io_enable_bits_taskID; // @[extracted_function_conv.scala 482:23]
  wire  const21_io_Out_ready; // @[extracted_function_conv.scala 482:23]
  wire  const21_io_Out_valid; // @[extracted_function_conv.scala 482:23]
  wire  const22_clock; // @[extracted_function_conv.scala 485:23]
  wire  const22_reset; // @[extracted_function_conv.scala 485:23]
  wire  const22_io_enable_ready; // @[extracted_function_conv.scala 485:23]
  wire  const22_io_enable_valid; // @[extracted_function_conv.scala 485:23]
  wire [4:0] const22_io_enable_bits_taskID; // @[extracted_function_conv.scala 485:23]
  wire  const22_io_Out_ready; // @[extracted_function_conv.scala 485:23]
  wire  const22_io_Out_valid; // @[extracted_function_conv.scala 485:23]
  wire  const23_clock; // @[extracted_function_conv.scala 488:23]
  wire  const23_reset; // @[extracted_function_conv.scala 488:23]
  wire  const23_io_enable_ready; // @[extracted_function_conv.scala 488:23]
  wire  const23_io_enable_valid; // @[extracted_function_conv.scala 488:23]
  wire [4:0] const23_io_enable_bits_taskID; // @[extracted_function_conv.scala 488:23]
  wire  const23_io_Out_ready; // @[extracted_function_conv.scala 488:23]
  wire  const23_io_Out_valid; // @[extracted_function_conv.scala 488:23]
  wire  const24_clock; // @[extracted_function_conv.scala 491:23]
  wire  const24_reset; // @[extracted_function_conv.scala 491:23]
  wire  const24_io_enable_ready; // @[extracted_function_conv.scala 491:23]
  wire  const24_io_enable_valid; // @[extracted_function_conv.scala 491:23]
  wire [4:0] const24_io_enable_bits_taskID; // @[extracted_function_conv.scala 491:23]
  wire  const24_io_Out_ready; // @[extracted_function_conv.scala 491:23]
  wire  const24_io_Out_valid; // @[extracted_function_conv.scala 491:23]
  wire  const25_clock; // @[extracted_function_conv.scala 494:23]
  wire  const25_reset; // @[extracted_function_conv.scala 494:23]
  wire  const25_io_enable_ready; // @[extracted_function_conv.scala 494:23]
  wire  const25_io_enable_valid; // @[extracted_function_conv.scala 494:23]
  wire [4:0] const25_io_enable_bits_taskID; // @[extracted_function_conv.scala 494:23]
  wire  const25_io_Out_ready; // @[extracted_function_conv.scala 494:23]
  wire  const25_io_Out_valid; // @[extracted_function_conv.scala 494:23]
  UnifiedController MemCtrl ( // @[extracted_function_conv.scala 45:23]
    .clock(MemCtrl_clock),
    .reset(MemCtrl_reset),
    .io_WriteIn_0_ready(MemCtrl_io_WriteIn_0_ready),
    .io_WriteIn_0_valid(MemCtrl_io_WriteIn_0_valid),
    .io_WriteIn_0_bits_address(MemCtrl_io_WriteIn_0_bits_address),
    .io_WriteIn_0_bits_data(MemCtrl_io_WriteIn_0_bits_data),
    .io_WriteIn_0_bits_taskID(MemCtrl_io_WriteIn_0_bits_taskID),
    .io_WriteIn_1_ready(MemCtrl_io_WriteIn_1_ready),
    .io_WriteIn_1_valid(MemCtrl_io_WriteIn_1_valid),
    .io_WriteIn_1_bits_address(MemCtrl_io_WriteIn_1_bits_address),
    .io_WriteIn_1_bits_data(MemCtrl_io_WriteIn_1_bits_data),
    .io_WriteIn_1_bits_taskID(MemCtrl_io_WriteIn_1_bits_taskID),
    .io_WriteIn_2_ready(MemCtrl_io_WriteIn_2_ready),
    .io_WriteIn_2_valid(MemCtrl_io_WriteIn_2_valid),
    .io_WriteIn_2_bits_address(MemCtrl_io_WriteIn_2_bits_address),
    .io_WriteIn_2_bits_data(MemCtrl_io_WriteIn_2_bits_data),
    .io_WriteIn_2_bits_taskID(MemCtrl_io_WriteIn_2_bits_taskID),
    .io_WriteIn_3_ready(MemCtrl_io_WriteIn_3_ready),
    .io_WriteIn_3_valid(MemCtrl_io_WriteIn_3_valid),
    .io_WriteIn_3_bits_address(MemCtrl_io_WriteIn_3_bits_address),
    .io_WriteIn_3_bits_data(MemCtrl_io_WriteIn_3_bits_data),
    .io_WriteIn_3_bits_taskID(MemCtrl_io_WriteIn_3_bits_taskID),
    .io_WriteIn_4_ready(MemCtrl_io_WriteIn_4_ready),
    .io_WriteIn_4_valid(MemCtrl_io_WriteIn_4_valid),
    .io_WriteIn_4_bits_address(MemCtrl_io_WriteIn_4_bits_address),
    .io_WriteIn_4_bits_data(MemCtrl_io_WriteIn_4_bits_data),
    .io_WriteIn_4_bits_taskID(MemCtrl_io_WriteIn_4_bits_taskID),
    .io_WriteIn_5_ready(MemCtrl_io_WriteIn_5_ready),
    .io_WriteIn_5_valid(MemCtrl_io_WriteIn_5_valid),
    .io_WriteIn_5_bits_address(MemCtrl_io_WriteIn_5_bits_address),
    .io_WriteIn_5_bits_data(MemCtrl_io_WriteIn_5_bits_data),
    .io_WriteIn_5_bits_taskID(MemCtrl_io_WriteIn_5_bits_taskID),
    .io_WriteIn_6_ready(MemCtrl_io_WriteIn_6_ready),
    .io_WriteIn_6_valid(MemCtrl_io_WriteIn_6_valid),
    .io_WriteIn_6_bits_address(MemCtrl_io_WriteIn_6_bits_address),
    .io_WriteIn_6_bits_data(MemCtrl_io_WriteIn_6_bits_data),
    .io_WriteIn_6_bits_taskID(MemCtrl_io_WriteIn_6_bits_taskID),
    .io_WriteIn_7_ready(MemCtrl_io_WriteIn_7_ready),
    .io_WriteIn_7_valid(MemCtrl_io_WriteIn_7_valid),
    .io_WriteIn_7_bits_address(MemCtrl_io_WriteIn_7_bits_address),
    .io_WriteIn_7_bits_data(MemCtrl_io_WriteIn_7_bits_data),
    .io_WriteIn_7_bits_taskID(MemCtrl_io_WriteIn_7_bits_taskID),
    .io_WriteIn_8_ready(MemCtrl_io_WriteIn_8_ready),
    .io_WriteIn_8_valid(MemCtrl_io_WriteIn_8_valid),
    .io_WriteIn_8_bits_address(MemCtrl_io_WriteIn_8_bits_address),
    .io_WriteIn_8_bits_data(MemCtrl_io_WriteIn_8_bits_data),
    .io_WriteIn_8_bits_taskID(MemCtrl_io_WriteIn_8_bits_taskID),
    .io_WriteOut_0_valid(MemCtrl_io_WriteOut_0_valid),
    .io_WriteOut_1_valid(MemCtrl_io_WriteOut_1_valid),
    .io_WriteOut_2_valid(MemCtrl_io_WriteOut_2_valid),
    .io_WriteOut_3_valid(MemCtrl_io_WriteOut_3_valid),
    .io_WriteOut_4_valid(MemCtrl_io_WriteOut_4_valid),
    .io_WriteOut_5_valid(MemCtrl_io_WriteOut_5_valid),
    .io_WriteOut_6_valid(MemCtrl_io_WriteOut_6_valid),
    .io_WriteOut_7_valid(MemCtrl_io_WriteOut_7_valid),
    .io_WriteOut_8_valid(MemCtrl_io_WriteOut_8_valid),
    .io_ReadIn_0_ready(MemCtrl_io_ReadIn_0_ready),
    .io_ReadIn_0_valid(MemCtrl_io_ReadIn_0_valid),
    .io_ReadIn_0_bits_address(MemCtrl_io_ReadIn_0_bits_address),
    .io_ReadIn_0_bits_taskID(MemCtrl_io_ReadIn_0_bits_taskID),
    .io_ReadIn_1_ready(MemCtrl_io_ReadIn_1_ready),
    .io_ReadIn_1_valid(MemCtrl_io_ReadIn_1_valid),
    .io_ReadIn_1_bits_address(MemCtrl_io_ReadIn_1_bits_address),
    .io_ReadIn_1_bits_taskID(MemCtrl_io_ReadIn_1_bits_taskID),
    .io_ReadIn_2_ready(MemCtrl_io_ReadIn_2_ready),
    .io_ReadIn_2_valid(MemCtrl_io_ReadIn_2_valid),
    .io_ReadIn_2_bits_address(MemCtrl_io_ReadIn_2_bits_address),
    .io_ReadIn_2_bits_taskID(MemCtrl_io_ReadIn_2_bits_taskID),
    .io_ReadIn_3_ready(MemCtrl_io_ReadIn_3_ready),
    .io_ReadIn_3_valid(MemCtrl_io_ReadIn_3_valid),
    .io_ReadIn_3_bits_address(MemCtrl_io_ReadIn_3_bits_address),
    .io_ReadIn_3_bits_taskID(MemCtrl_io_ReadIn_3_bits_taskID),
    .io_ReadIn_4_ready(MemCtrl_io_ReadIn_4_ready),
    .io_ReadIn_4_valid(MemCtrl_io_ReadIn_4_valid),
    .io_ReadIn_4_bits_address(MemCtrl_io_ReadIn_4_bits_address),
    .io_ReadIn_4_bits_taskID(MemCtrl_io_ReadIn_4_bits_taskID),
    .io_ReadIn_5_ready(MemCtrl_io_ReadIn_5_ready),
    .io_ReadIn_5_valid(MemCtrl_io_ReadIn_5_valid),
    .io_ReadIn_5_bits_address(MemCtrl_io_ReadIn_5_bits_address),
    .io_ReadIn_5_bits_taskID(MemCtrl_io_ReadIn_5_bits_taskID),
    .io_ReadIn_6_ready(MemCtrl_io_ReadIn_6_ready),
    .io_ReadIn_6_valid(MemCtrl_io_ReadIn_6_valid),
    .io_ReadIn_6_bits_address(MemCtrl_io_ReadIn_6_bits_address),
    .io_ReadIn_6_bits_taskID(MemCtrl_io_ReadIn_6_bits_taskID),
    .io_ReadIn_7_ready(MemCtrl_io_ReadIn_7_ready),
    .io_ReadIn_7_valid(MemCtrl_io_ReadIn_7_valid),
    .io_ReadIn_7_bits_address(MemCtrl_io_ReadIn_7_bits_address),
    .io_ReadIn_7_bits_taskID(MemCtrl_io_ReadIn_7_bits_taskID),
    .io_ReadIn_8_ready(MemCtrl_io_ReadIn_8_ready),
    .io_ReadIn_8_valid(MemCtrl_io_ReadIn_8_valid),
    .io_ReadIn_8_bits_address(MemCtrl_io_ReadIn_8_bits_address),
    .io_ReadIn_8_bits_taskID(MemCtrl_io_ReadIn_8_bits_taskID),
    .io_ReadIn_9_ready(MemCtrl_io_ReadIn_9_ready),
    .io_ReadIn_9_valid(MemCtrl_io_ReadIn_9_valid),
    .io_ReadIn_9_bits_address(MemCtrl_io_ReadIn_9_bits_address),
    .io_ReadIn_9_bits_taskID(MemCtrl_io_ReadIn_9_bits_taskID),
    .io_ReadIn_10_ready(MemCtrl_io_ReadIn_10_ready),
    .io_ReadIn_10_valid(MemCtrl_io_ReadIn_10_valid),
    .io_ReadIn_10_bits_address(MemCtrl_io_ReadIn_10_bits_address),
    .io_ReadIn_10_bits_taskID(MemCtrl_io_ReadIn_10_bits_taskID),
    .io_ReadIn_11_ready(MemCtrl_io_ReadIn_11_ready),
    .io_ReadIn_11_valid(MemCtrl_io_ReadIn_11_valid),
    .io_ReadIn_11_bits_address(MemCtrl_io_ReadIn_11_bits_address),
    .io_ReadIn_11_bits_taskID(MemCtrl_io_ReadIn_11_bits_taskID),
    .io_ReadIn_12_ready(MemCtrl_io_ReadIn_12_ready),
    .io_ReadIn_12_valid(MemCtrl_io_ReadIn_12_valid),
    .io_ReadIn_12_bits_address(MemCtrl_io_ReadIn_12_bits_address),
    .io_ReadIn_12_bits_taskID(MemCtrl_io_ReadIn_12_bits_taskID),
    .io_ReadIn_13_ready(MemCtrl_io_ReadIn_13_ready),
    .io_ReadIn_13_valid(MemCtrl_io_ReadIn_13_valid),
    .io_ReadIn_13_bits_address(MemCtrl_io_ReadIn_13_bits_address),
    .io_ReadIn_13_bits_taskID(MemCtrl_io_ReadIn_13_bits_taskID),
    .io_ReadIn_14_ready(MemCtrl_io_ReadIn_14_ready),
    .io_ReadIn_14_valid(MemCtrl_io_ReadIn_14_valid),
    .io_ReadIn_14_bits_address(MemCtrl_io_ReadIn_14_bits_address),
    .io_ReadIn_14_bits_taskID(MemCtrl_io_ReadIn_14_bits_taskID),
    .io_ReadIn_15_ready(MemCtrl_io_ReadIn_15_ready),
    .io_ReadIn_15_valid(MemCtrl_io_ReadIn_15_valid),
    .io_ReadIn_15_bits_address(MemCtrl_io_ReadIn_15_bits_address),
    .io_ReadIn_15_bits_taskID(MemCtrl_io_ReadIn_15_bits_taskID),
    .io_ReadIn_16_ready(MemCtrl_io_ReadIn_16_ready),
    .io_ReadIn_16_valid(MemCtrl_io_ReadIn_16_valid),
    .io_ReadIn_16_bits_address(MemCtrl_io_ReadIn_16_bits_address),
    .io_ReadIn_16_bits_taskID(MemCtrl_io_ReadIn_16_bits_taskID),
    .io_ReadIn_17_ready(MemCtrl_io_ReadIn_17_ready),
    .io_ReadIn_17_valid(MemCtrl_io_ReadIn_17_valid),
    .io_ReadIn_17_bits_address(MemCtrl_io_ReadIn_17_bits_address),
    .io_ReadIn_17_bits_taskID(MemCtrl_io_ReadIn_17_bits_taskID),
    .io_ReadIn_18_ready(MemCtrl_io_ReadIn_18_ready),
    .io_ReadIn_18_valid(MemCtrl_io_ReadIn_18_valid),
    .io_ReadIn_18_bits_address(MemCtrl_io_ReadIn_18_bits_address),
    .io_ReadIn_18_bits_taskID(MemCtrl_io_ReadIn_18_bits_taskID),
    .io_ReadOut_0_valid(MemCtrl_io_ReadOut_0_valid),
    .io_ReadOut_0_data(MemCtrl_io_ReadOut_0_data),
    .io_ReadOut_1_valid(MemCtrl_io_ReadOut_1_valid),
    .io_ReadOut_1_data(MemCtrl_io_ReadOut_1_data),
    .io_ReadOut_2_valid(MemCtrl_io_ReadOut_2_valid),
    .io_ReadOut_2_data(MemCtrl_io_ReadOut_2_data),
    .io_ReadOut_3_valid(MemCtrl_io_ReadOut_3_valid),
    .io_ReadOut_3_data(MemCtrl_io_ReadOut_3_data),
    .io_ReadOut_4_valid(MemCtrl_io_ReadOut_4_valid),
    .io_ReadOut_4_data(MemCtrl_io_ReadOut_4_data),
    .io_ReadOut_5_valid(MemCtrl_io_ReadOut_5_valid),
    .io_ReadOut_5_data(MemCtrl_io_ReadOut_5_data),
    .io_ReadOut_6_valid(MemCtrl_io_ReadOut_6_valid),
    .io_ReadOut_6_data(MemCtrl_io_ReadOut_6_data),
    .io_ReadOut_7_valid(MemCtrl_io_ReadOut_7_valid),
    .io_ReadOut_7_data(MemCtrl_io_ReadOut_7_data),
    .io_ReadOut_8_valid(MemCtrl_io_ReadOut_8_valid),
    .io_ReadOut_8_data(MemCtrl_io_ReadOut_8_data),
    .io_ReadOut_9_valid(MemCtrl_io_ReadOut_9_valid),
    .io_ReadOut_9_data(MemCtrl_io_ReadOut_9_data),
    .io_ReadOut_10_valid(MemCtrl_io_ReadOut_10_valid),
    .io_ReadOut_10_data(MemCtrl_io_ReadOut_10_data),
    .io_ReadOut_11_valid(MemCtrl_io_ReadOut_11_valid),
    .io_ReadOut_11_data(MemCtrl_io_ReadOut_11_data),
    .io_ReadOut_12_valid(MemCtrl_io_ReadOut_12_valid),
    .io_ReadOut_12_data(MemCtrl_io_ReadOut_12_data),
    .io_ReadOut_13_valid(MemCtrl_io_ReadOut_13_valid),
    .io_ReadOut_13_data(MemCtrl_io_ReadOut_13_data),
    .io_ReadOut_14_valid(MemCtrl_io_ReadOut_14_valid),
    .io_ReadOut_14_data(MemCtrl_io_ReadOut_14_data),
    .io_ReadOut_15_valid(MemCtrl_io_ReadOut_15_valid),
    .io_ReadOut_15_data(MemCtrl_io_ReadOut_15_data),
    .io_ReadOut_16_valid(MemCtrl_io_ReadOut_16_valid),
    .io_ReadOut_16_data(MemCtrl_io_ReadOut_16_data),
    .io_ReadOut_17_valid(MemCtrl_io_ReadOut_17_valid),
    .io_ReadOut_17_data(MemCtrl_io_ReadOut_17_data),
    .io_ReadOut_18_valid(MemCtrl_io_ReadOut_18_valid),
    .io_ReadOut_18_data(MemCtrl_io_ReadOut_18_data),
    .io_MemResp_valid(MemCtrl_io_MemResp_valid),
    .io_MemResp_bits_data(MemCtrl_io_MemResp_bits_data),
    .io_MemResp_bits_tag(MemCtrl_io_MemResp_bits_tag),
    .io_MemResp_bits_iswrite(MemCtrl_io_MemResp_bits_iswrite),
    .io_MemReq_ready(MemCtrl_io_MemReq_ready),
    .io_MemReq_valid(MemCtrl_io_MemReq_valid),
    .io_MemReq_bits_addr(MemCtrl_io_MemReq_bits_addr),
    .io_MemReq_bits_data(MemCtrl_io_MemReq_bits_data),
    .io_MemReq_bits_mask(MemCtrl_io_MemReq_bits_mask),
    .io_MemReq_bits_tag(MemCtrl_io_MemReq_bits_tag),
    .io_MemReq_bits_taskID(MemCtrl_io_MemReq_bits_taskID),
    .io_MemReq_bits_iswrite(MemCtrl_io_MemReq_bits_iswrite)
  );
  SplitCallNew InputSplitter ( // @[extracted_function_conv.scala 53:29]
    .clock(InputSplitter_clock),
    .reset(InputSplitter_reset),
    .io_In_ready(InputSplitter_io_In_ready),
    .io_In_valid(InputSplitter_io_In_valid),
    .io_In_bits_enable_taskID(InputSplitter_io_In_bits_enable_taskID),
    .io_In_bits_enable_control(InputSplitter_io_In_bits_enable_control),
    .io_In_bits_data_field5_data(InputSplitter_io_In_bits_data_field5_data),
    .io_In_bits_data_field4_data(InputSplitter_io_In_bits_data_field4_data),
    .io_In_bits_data_field3_data(InputSplitter_io_In_bits_data_field3_data),
    .io_In_bits_data_field2_taskID(InputSplitter_io_In_bits_data_field2_taskID),
    .io_In_bits_data_field2_data(InputSplitter_io_In_bits_data_field2_data),
    .io_In_bits_data_field1_predicate(InputSplitter_io_In_bits_data_field1_predicate),
    .io_In_bits_data_field1_taskID(InputSplitter_io_In_bits_data_field1_taskID),
    .io_In_bits_data_field1_data(InputSplitter_io_In_bits_data_field1_data),
    .io_In_bits_data_field0_taskID(InputSplitter_io_In_bits_data_field0_taskID),
    .io_In_bits_data_field0_data(InputSplitter_io_In_bits_data_field0_data),
    .io_Out_enable_ready(InputSplitter_io_Out_enable_ready),
    .io_Out_enable_valid(InputSplitter_io_Out_enable_valid),
    .io_Out_enable_bits_taskID(InputSplitter_io_Out_enable_bits_taskID),
    .io_Out_enable_bits_control(InputSplitter_io_Out_enable_bits_control),
    .io_Out_data_field5_0_ready(InputSplitter_io_Out_data_field5_0_ready),
    .io_Out_data_field5_0_valid(InputSplitter_io_Out_data_field5_0_valid),
    .io_Out_data_field5_0_bits_data(InputSplitter_io_Out_data_field5_0_bits_data),
    .io_Out_data_field5_1_ready(InputSplitter_io_Out_data_field5_1_ready),
    .io_Out_data_field5_1_valid(InputSplitter_io_Out_data_field5_1_valid),
    .io_Out_data_field5_1_bits_data(InputSplitter_io_Out_data_field5_1_bits_data),
    .io_Out_data_field4_0_ready(InputSplitter_io_Out_data_field4_0_ready),
    .io_Out_data_field4_0_valid(InputSplitter_io_Out_data_field4_0_valid),
    .io_Out_data_field4_0_bits_data(InputSplitter_io_Out_data_field4_0_bits_data),
    .io_Out_data_field3_0_ready(InputSplitter_io_Out_data_field3_0_ready),
    .io_Out_data_field3_0_valid(InputSplitter_io_Out_data_field3_0_valid),
    .io_Out_data_field3_0_bits_data(InputSplitter_io_Out_data_field3_0_bits_data),
    .io_Out_data_field2_0_ready(InputSplitter_io_Out_data_field2_0_ready),
    .io_Out_data_field2_0_valid(InputSplitter_io_Out_data_field2_0_valid),
    .io_Out_data_field2_0_bits_taskID(InputSplitter_io_Out_data_field2_0_bits_taskID),
    .io_Out_data_field2_0_bits_data(InputSplitter_io_Out_data_field2_0_bits_data),
    .io_Out_data_field1_0_ready(InputSplitter_io_Out_data_field1_0_ready),
    .io_Out_data_field1_0_valid(InputSplitter_io_Out_data_field1_0_valid),
    .io_Out_data_field1_0_bits_predicate(InputSplitter_io_Out_data_field1_0_bits_predicate),
    .io_Out_data_field1_0_bits_taskID(InputSplitter_io_Out_data_field1_0_bits_taskID),
    .io_Out_data_field1_0_bits_data(InputSplitter_io_Out_data_field1_0_bits_data),
    .io_Out_data_field1_1_ready(InputSplitter_io_Out_data_field1_1_ready),
    .io_Out_data_field1_1_valid(InputSplitter_io_Out_data_field1_1_valid),
    .io_Out_data_field1_1_bits_taskID(InputSplitter_io_Out_data_field1_1_bits_taskID),
    .io_Out_data_field1_1_bits_data(InputSplitter_io_Out_data_field1_1_bits_data),
    .io_Out_data_field1_2_ready(InputSplitter_io_Out_data_field1_2_ready),
    .io_Out_data_field1_2_valid(InputSplitter_io_Out_data_field1_2_valid),
    .io_Out_data_field1_2_bits_taskID(InputSplitter_io_Out_data_field1_2_bits_taskID),
    .io_Out_data_field1_2_bits_data(InputSplitter_io_Out_data_field1_2_bits_data),
    .io_Out_data_field1_3_ready(InputSplitter_io_Out_data_field1_3_ready),
    .io_Out_data_field1_3_valid(InputSplitter_io_Out_data_field1_3_valid),
    .io_Out_data_field1_3_bits_taskID(InputSplitter_io_Out_data_field1_3_bits_taskID),
    .io_Out_data_field1_3_bits_data(InputSplitter_io_Out_data_field1_3_bits_data),
    .io_Out_data_field1_4_ready(InputSplitter_io_Out_data_field1_4_ready),
    .io_Out_data_field1_4_valid(InputSplitter_io_Out_data_field1_4_valid),
    .io_Out_data_field1_4_bits_taskID(InputSplitter_io_Out_data_field1_4_bits_taskID),
    .io_Out_data_field1_4_bits_data(InputSplitter_io_Out_data_field1_4_bits_data),
    .io_Out_data_field1_5_ready(InputSplitter_io_Out_data_field1_5_ready),
    .io_Out_data_field1_5_valid(InputSplitter_io_Out_data_field1_5_valid),
    .io_Out_data_field1_5_bits_taskID(InputSplitter_io_Out_data_field1_5_bits_taskID),
    .io_Out_data_field1_5_bits_data(InputSplitter_io_Out_data_field1_5_bits_data),
    .io_Out_data_field1_6_ready(InputSplitter_io_Out_data_field1_6_ready),
    .io_Out_data_field1_6_valid(InputSplitter_io_Out_data_field1_6_valid),
    .io_Out_data_field1_6_bits_taskID(InputSplitter_io_Out_data_field1_6_bits_taskID),
    .io_Out_data_field1_6_bits_data(InputSplitter_io_Out_data_field1_6_bits_data),
    .io_Out_data_field1_7_ready(InputSplitter_io_Out_data_field1_7_ready),
    .io_Out_data_field1_7_valid(InputSplitter_io_Out_data_field1_7_valid),
    .io_Out_data_field1_7_bits_taskID(InputSplitter_io_Out_data_field1_7_bits_taskID),
    .io_Out_data_field1_7_bits_data(InputSplitter_io_Out_data_field1_7_bits_data),
    .io_Out_data_field1_8_ready(InputSplitter_io_Out_data_field1_8_ready),
    .io_Out_data_field1_8_valid(InputSplitter_io_Out_data_field1_8_valid),
    .io_Out_data_field1_8_bits_taskID(InputSplitter_io_Out_data_field1_8_bits_taskID),
    .io_Out_data_field1_8_bits_data(InputSplitter_io_Out_data_field1_8_bits_data),
    .io_Out_data_field0_0_ready(InputSplitter_io_Out_data_field0_0_ready),
    .io_Out_data_field0_0_valid(InputSplitter_io_Out_data_field0_0_valid),
    .io_Out_data_field0_0_bits_taskID(InputSplitter_io_Out_data_field0_0_bits_taskID),
    .io_Out_data_field0_0_bits_data(InputSplitter_io_Out_data_field0_0_bits_data)
  );
  LoopBlockNode Loop_0 ( // @[extracted_function_conv.scala 62:22]
    .clock(Loop_0_clock),
    .reset(Loop_0_reset),
    .io_enable_ready(Loop_0_io_enable_ready),
    .io_enable_valid(Loop_0_io_enable_valid),
    .io_enable_bits_taskID(Loop_0_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_0_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_0_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_0_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_0_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_0_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_0_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_0_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_0_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_0_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_data(Loop_0_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_0_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_0_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_data(Loop_0_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_0_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_0_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_predicate(Loop_0_io_InLiveIn_4_bits_predicate),
    .io_InLiveIn_4_bits_taskID(Loop_0_io_InLiveIn_4_bits_taskID),
    .io_InLiveIn_4_bits_data(Loop_0_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_0_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_0_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_data(Loop_0_io_InLiveIn_5_bits_data),
    .io_InLiveIn_6_ready(Loop_0_io_InLiveIn_6_ready),
    .io_InLiveIn_6_valid(Loop_0_io_InLiveIn_6_valid),
    .io_InLiveIn_6_bits_predicate(Loop_0_io_InLiveIn_6_bits_predicate),
    .io_InLiveIn_6_bits_taskID(Loop_0_io_InLiveIn_6_bits_taskID),
    .io_InLiveIn_6_bits_data(Loop_0_io_InLiveIn_6_bits_data),
    .io_InLiveIn_7_ready(Loop_0_io_InLiveIn_7_ready),
    .io_InLiveIn_7_valid(Loop_0_io_InLiveIn_7_valid),
    .io_InLiveIn_7_bits_predicate(Loop_0_io_InLiveIn_7_bits_predicate),
    .io_InLiveIn_7_bits_taskID(Loop_0_io_InLiveIn_7_bits_taskID),
    .io_InLiveIn_7_bits_data(Loop_0_io_InLiveIn_7_bits_data),
    .io_InLiveIn_8_ready(Loop_0_io_InLiveIn_8_ready),
    .io_InLiveIn_8_valid(Loop_0_io_InLiveIn_8_valid),
    .io_InLiveIn_8_bits_predicate(Loop_0_io_InLiveIn_8_bits_predicate),
    .io_InLiveIn_8_bits_taskID(Loop_0_io_InLiveIn_8_bits_taskID),
    .io_InLiveIn_8_bits_data(Loop_0_io_InLiveIn_8_bits_data),
    .io_InLiveIn_9_ready(Loop_0_io_InLiveIn_9_ready),
    .io_InLiveIn_9_valid(Loop_0_io_InLiveIn_9_valid),
    .io_InLiveIn_9_bits_predicate(Loop_0_io_InLiveIn_9_bits_predicate),
    .io_InLiveIn_9_bits_taskID(Loop_0_io_InLiveIn_9_bits_taskID),
    .io_InLiveIn_9_bits_data(Loop_0_io_InLiveIn_9_bits_data),
    .io_InLiveIn_10_ready(Loop_0_io_InLiveIn_10_ready),
    .io_InLiveIn_10_valid(Loop_0_io_InLiveIn_10_valid),
    .io_InLiveIn_10_bits_taskID(Loop_0_io_InLiveIn_10_bits_taskID),
    .io_InLiveIn_10_bits_data(Loop_0_io_InLiveIn_10_bits_data),
    .io_InLiveIn_11_ready(Loop_0_io_InLiveIn_11_ready),
    .io_InLiveIn_11_valid(Loop_0_io_InLiveIn_11_valid),
    .io_InLiveIn_11_bits_taskID(Loop_0_io_InLiveIn_11_bits_taskID),
    .io_InLiveIn_11_bits_data(Loop_0_io_InLiveIn_11_bits_data),
    .io_InLiveIn_12_ready(Loop_0_io_InLiveIn_12_ready),
    .io_InLiveIn_12_valid(Loop_0_io_InLiveIn_12_valid),
    .io_InLiveIn_12_bits_predicate(Loop_0_io_InLiveIn_12_bits_predicate),
    .io_InLiveIn_12_bits_taskID(Loop_0_io_InLiveIn_12_bits_taskID),
    .io_InLiveIn_12_bits_data(Loop_0_io_InLiveIn_12_bits_data),
    .io_InLiveIn_13_ready(Loop_0_io_InLiveIn_13_ready),
    .io_InLiveIn_13_valid(Loop_0_io_InLiveIn_13_valid),
    .io_InLiveIn_13_bits_predicate(Loop_0_io_InLiveIn_13_bits_predicate),
    .io_InLiveIn_13_bits_taskID(Loop_0_io_InLiveIn_13_bits_taskID),
    .io_InLiveIn_13_bits_data(Loop_0_io_InLiveIn_13_bits_data),
    .io_InLiveIn_14_ready(Loop_0_io_InLiveIn_14_ready),
    .io_InLiveIn_14_valid(Loop_0_io_InLiveIn_14_valid),
    .io_InLiveIn_14_bits_predicate(Loop_0_io_InLiveIn_14_bits_predicate),
    .io_InLiveIn_14_bits_taskID(Loop_0_io_InLiveIn_14_bits_taskID),
    .io_InLiveIn_14_bits_data(Loop_0_io_InLiveIn_14_bits_data),
    .io_InLiveIn_15_ready(Loop_0_io_InLiveIn_15_ready),
    .io_InLiveIn_15_valid(Loop_0_io_InLiveIn_15_valid),
    .io_InLiveIn_15_bits_predicate(Loop_0_io_InLiveIn_15_bits_predicate),
    .io_InLiveIn_15_bits_taskID(Loop_0_io_InLiveIn_15_bits_taskID),
    .io_InLiveIn_15_bits_data(Loop_0_io_InLiveIn_15_bits_data),
    .io_OutLiveIn_field15_0_ready(Loop_0_io_OutLiveIn_field15_0_ready),
    .io_OutLiveIn_field15_0_valid(Loop_0_io_OutLiveIn_field15_0_valid),
    .io_OutLiveIn_field15_0_bits_predicate(Loop_0_io_OutLiveIn_field15_0_bits_predicate),
    .io_OutLiveIn_field15_0_bits_taskID(Loop_0_io_OutLiveIn_field15_0_bits_taskID),
    .io_OutLiveIn_field15_0_bits_data(Loop_0_io_OutLiveIn_field15_0_bits_data),
    .io_OutLiveIn_field14_0_ready(Loop_0_io_OutLiveIn_field14_0_ready),
    .io_OutLiveIn_field14_0_valid(Loop_0_io_OutLiveIn_field14_0_valid),
    .io_OutLiveIn_field14_0_bits_predicate(Loop_0_io_OutLiveIn_field14_0_bits_predicate),
    .io_OutLiveIn_field14_0_bits_taskID(Loop_0_io_OutLiveIn_field14_0_bits_taskID),
    .io_OutLiveIn_field14_0_bits_data(Loop_0_io_OutLiveIn_field14_0_bits_data),
    .io_OutLiveIn_field13_0_ready(Loop_0_io_OutLiveIn_field13_0_ready),
    .io_OutLiveIn_field13_0_valid(Loop_0_io_OutLiveIn_field13_0_valid),
    .io_OutLiveIn_field13_0_bits_predicate(Loop_0_io_OutLiveIn_field13_0_bits_predicate),
    .io_OutLiveIn_field13_0_bits_taskID(Loop_0_io_OutLiveIn_field13_0_bits_taskID),
    .io_OutLiveIn_field13_0_bits_data(Loop_0_io_OutLiveIn_field13_0_bits_data),
    .io_OutLiveIn_field12_0_ready(Loop_0_io_OutLiveIn_field12_0_ready),
    .io_OutLiveIn_field12_0_valid(Loop_0_io_OutLiveIn_field12_0_valid),
    .io_OutLiveIn_field12_0_bits_predicate(Loop_0_io_OutLiveIn_field12_0_bits_predicate),
    .io_OutLiveIn_field12_0_bits_taskID(Loop_0_io_OutLiveIn_field12_0_bits_taskID),
    .io_OutLiveIn_field12_0_bits_data(Loop_0_io_OutLiveIn_field12_0_bits_data),
    .io_OutLiveIn_field11_0_ready(Loop_0_io_OutLiveIn_field11_0_ready),
    .io_OutLiveIn_field11_0_valid(Loop_0_io_OutLiveIn_field11_0_valid),
    .io_OutLiveIn_field11_0_bits_taskID(Loop_0_io_OutLiveIn_field11_0_bits_taskID),
    .io_OutLiveIn_field11_0_bits_data(Loop_0_io_OutLiveIn_field11_0_bits_data),
    .io_OutLiveIn_field10_0_ready(Loop_0_io_OutLiveIn_field10_0_ready),
    .io_OutLiveIn_field10_0_valid(Loop_0_io_OutLiveIn_field10_0_valid),
    .io_OutLiveIn_field10_0_bits_taskID(Loop_0_io_OutLiveIn_field10_0_bits_taskID),
    .io_OutLiveIn_field10_0_bits_data(Loop_0_io_OutLiveIn_field10_0_bits_data),
    .io_OutLiveIn_field10_1_ready(Loop_0_io_OutLiveIn_field10_1_ready),
    .io_OutLiveIn_field10_1_valid(Loop_0_io_OutLiveIn_field10_1_valid),
    .io_OutLiveIn_field10_1_bits_taskID(Loop_0_io_OutLiveIn_field10_1_bits_taskID),
    .io_OutLiveIn_field10_1_bits_data(Loop_0_io_OutLiveIn_field10_1_bits_data),
    .io_OutLiveIn_field10_2_ready(Loop_0_io_OutLiveIn_field10_2_ready),
    .io_OutLiveIn_field10_2_valid(Loop_0_io_OutLiveIn_field10_2_valid),
    .io_OutLiveIn_field10_2_bits_taskID(Loop_0_io_OutLiveIn_field10_2_bits_taskID),
    .io_OutLiveIn_field10_2_bits_data(Loop_0_io_OutLiveIn_field10_2_bits_data),
    .io_OutLiveIn_field10_3_ready(Loop_0_io_OutLiveIn_field10_3_ready),
    .io_OutLiveIn_field10_3_valid(Loop_0_io_OutLiveIn_field10_3_valid),
    .io_OutLiveIn_field10_3_bits_taskID(Loop_0_io_OutLiveIn_field10_3_bits_taskID),
    .io_OutLiveIn_field10_3_bits_data(Loop_0_io_OutLiveIn_field10_3_bits_data),
    .io_OutLiveIn_field10_4_ready(Loop_0_io_OutLiveIn_field10_4_ready),
    .io_OutLiveIn_field10_4_valid(Loop_0_io_OutLiveIn_field10_4_valid),
    .io_OutLiveIn_field10_4_bits_taskID(Loop_0_io_OutLiveIn_field10_4_bits_taskID),
    .io_OutLiveIn_field10_4_bits_data(Loop_0_io_OutLiveIn_field10_4_bits_data),
    .io_OutLiveIn_field10_5_ready(Loop_0_io_OutLiveIn_field10_5_ready),
    .io_OutLiveIn_field10_5_valid(Loop_0_io_OutLiveIn_field10_5_valid),
    .io_OutLiveIn_field10_5_bits_taskID(Loop_0_io_OutLiveIn_field10_5_bits_taskID),
    .io_OutLiveIn_field10_5_bits_data(Loop_0_io_OutLiveIn_field10_5_bits_data),
    .io_OutLiveIn_field10_6_ready(Loop_0_io_OutLiveIn_field10_6_ready),
    .io_OutLiveIn_field10_6_valid(Loop_0_io_OutLiveIn_field10_6_valid),
    .io_OutLiveIn_field10_6_bits_taskID(Loop_0_io_OutLiveIn_field10_6_bits_taskID),
    .io_OutLiveIn_field10_6_bits_data(Loop_0_io_OutLiveIn_field10_6_bits_data),
    .io_OutLiveIn_field10_7_ready(Loop_0_io_OutLiveIn_field10_7_ready),
    .io_OutLiveIn_field10_7_valid(Loop_0_io_OutLiveIn_field10_7_valid),
    .io_OutLiveIn_field10_7_bits_taskID(Loop_0_io_OutLiveIn_field10_7_bits_taskID),
    .io_OutLiveIn_field10_7_bits_data(Loop_0_io_OutLiveIn_field10_7_bits_data),
    .io_OutLiveIn_field10_8_ready(Loop_0_io_OutLiveIn_field10_8_ready),
    .io_OutLiveIn_field10_8_valid(Loop_0_io_OutLiveIn_field10_8_valid),
    .io_OutLiveIn_field10_8_bits_taskID(Loop_0_io_OutLiveIn_field10_8_bits_taskID),
    .io_OutLiveIn_field10_8_bits_data(Loop_0_io_OutLiveIn_field10_8_bits_data),
    .io_OutLiveIn_field9_0_ready(Loop_0_io_OutLiveIn_field9_0_ready),
    .io_OutLiveIn_field9_0_valid(Loop_0_io_OutLiveIn_field9_0_valid),
    .io_OutLiveIn_field9_0_bits_predicate(Loop_0_io_OutLiveIn_field9_0_bits_predicate),
    .io_OutLiveIn_field9_0_bits_taskID(Loop_0_io_OutLiveIn_field9_0_bits_taskID),
    .io_OutLiveIn_field9_0_bits_data(Loop_0_io_OutLiveIn_field9_0_bits_data),
    .io_OutLiveIn_field8_0_ready(Loop_0_io_OutLiveIn_field8_0_ready),
    .io_OutLiveIn_field8_0_valid(Loop_0_io_OutLiveIn_field8_0_valid),
    .io_OutLiveIn_field8_0_bits_predicate(Loop_0_io_OutLiveIn_field8_0_bits_predicate),
    .io_OutLiveIn_field8_0_bits_taskID(Loop_0_io_OutLiveIn_field8_0_bits_taskID),
    .io_OutLiveIn_field8_0_bits_data(Loop_0_io_OutLiveIn_field8_0_bits_data),
    .io_OutLiveIn_field7_0_ready(Loop_0_io_OutLiveIn_field7_0_ready),
    .io_OutLiveIn_field7_0_valid(Loop_0_io_OutLiveIn_field7_0_valid),
    .io_OutLiveIn_field7_0_bits_predicate(Loop_0_io_OutLiveIn_field7_0_bits_predicate),
    .io_OutLiveIn_field7_0_bits_taskID(Loop_0_io_OutLiveIn_field7_0_bits_taskID),
    .io_OutLiveIn_field7_0_bits_data(Loop_0_io_OutLiveIn_field7_0_bits_data),
    .io_OutLiveIn_field6_0_ready(Loop_0_io_OutLiveIn_field6_0_ready),
    .io_OutLiveIn_field6_0_valid(Loop_0_io_OutLiveIn_field6_0_valid),
    .io_OutLiveIn_field6_0_bits_predicate(Loop_0_io_OutLiveIn_field6_0_bits_predicate),
    .io_OutLiveIn_field6_0_bits_taskID(Loop_0_io_OutLiveIn_field6_0_bits_taskID),
    .io_OutLiveIn_field6_0_bits_data(Loop_0_io_OutLiveIn_field6_0_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_0_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_0_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_data(Loop_0_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_0_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_0_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_predicate(Loop_0_io_OutLiveIn_field4_0_bits_predicate),
    .io_OutLiveIn_field4_0_bits_taskID(Loop_0_io_OutLiveIn_field4_0_bits_taskID),
    .io_OutLiveIn_field4_0_bits_data(Loop_0_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_0_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_0_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_data(Loop_0_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_0_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_0_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_data(Loop_0_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_0_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_0_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_0_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_0_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_0_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_0_io_OutLiveIn_field0_0_bits_data),
    .io_activate_loop_start_ready(Loop_0_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_0_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_0_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_0_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_0_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_0_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_0_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_0_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_0_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_0_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_0_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_0_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_0_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_0_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_0_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_0_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_0_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_0_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_0_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_0_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_0_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_0_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_0_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_0_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_0_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_0_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_0_io_loopExit_0_bits_control)
  );
  LoopBlockNode_1 Loop_1 ( // @[extracted_function_conv.scala 64:22]
    .clock(Loop_1_clock),
    .reset(Loop_1_reset),
    .io_enable_ready(Loop_1_io_enable_ready),
    .io_enable_valid(Loop_1_io_enable_valid),
    .io_enable_bits_taskID(Loop_1_io_enable_bits_taskID),
    .io_enable_bits_control(Loop_1_io_enable_bits_control),
    .io_InLiveIn_0_ready(Loop_1_io_InLiveIn_0_ready),
    .io_InLiveIn_0_valid(Loop_1_io_InLiveIn_0_valid),
    .io_InLiveIn_0_bits_data(Loop_1_io_InLiveIn_0_bits_data),
    .io_InLiveIn_1_ready(Loop_1_io_InLiveIn_1_ready),
    .io_InLiveIn_1_valid(Loop_1_io_InLiveIn_1_valid),
    .io_InLiveIn_1_bits_data(Loop_1_io_InLiveIn_1_bits_data),
    .io_InLiveIn_2_ready(Loop_1_io_InLiveIn_2_ready),
    .io_InLiveIn_2_valid(Loop_1_io_InLiveIn_2_valid),
    .io_InLiveIn_2_bits_taskID(Loop_1_io_InLiveIn_2_bits_taskID),
    .io_InLiveIn_2_bits_data(Loop_1_io_InLiveIn_2_bits_data),
    .io_InLiveIn_3_ready(Loop_1_io_InLiveIn_3_ready),
    .io_InLiveIn_3_valid(Loop_1_io_InLiveIn_3_valid),
    .io_InLiveIn_3_bits_predicate(Loop_1_io_InLiveIn_3_bits_predicate),
    .io_InLiveIn_3_bits_taskID(Loop_1_io_InLiveIn_3_bits_taskID),
    .io_InLiveIn_3_bits_data(Loop_1_io_InLiveIn_3_bits_data),
    .io_InLiveIn_4_ready(Loop_1_io_InLiveIn_4_ready),
    .io_InLiveIn_4_valid(Loop_1_io_InLiveIn_4_valid),
    .io_InLiveIn_4_bits_taskID(Loop_1_io_InLiveIn_4_bits_taskID),
    .io_InLiveIn_4_bits_data(Loop_1_io_InLiveIn_4_bits_data),
    .io_InLiveIn_5_ready(Loop_1_io_InLiveIn_5_ready),
    .io_InLiveIn_5_valid(Loop_1_io_InLiveIn_5_valid),
    .io_InLiveIn_5_bits_predicate(Loop_1_io_InLiveIn_5_bits_predicate),
    .io_InLiveIn_5_bits_taskID(Loop_1_io_InLiveIn_5_bits_taskID),
    .io_InLiveIn_5_bits_data(Loop_1_io_InLiveIn_5_bits_data),
    .io_InLiveIn_6_ready(Loop_1_io_InLiveIn_6_ready),
    .io_InLiveIn_6_valid(Loop_1_io_InLiveIn_6_valid),
    .io_InLiveIn_6_bits_predicate(Loop_1_io_InLiveIn_6_bits_predicate),
    .io_InLiveIn_6_bits_taskID(Loop_1_io_InLiveIn_6_bits_taskID),
    .io_InLiveIn_6_bits_data(Loop_1_io_InLiveIn_6_bits_data),
    .io_InLiveIn_7_ready(Loop_1_io_InLiveIn_7_ready),
    .io_InLiveIn_7_valid(Loop_1_io_InLiveIn_7_valid),
    .io_InLiveIn_7_bits_predicate(Loop_1_io_InLiveIn_7_bits_predicate),
    .io_InLiveIn_7_bits_taskID(Loop_1_io_InLiveIn_7_bits_taskID),
    .io_InLiveIn_7_bits_data(Loop_1_io_InLiveIn_7_bits_data),
    .io_InLiveIn_8_ready(Loop_1_io_InLiveIn_8_ready),
    .io_InLiveIn_8_valid(Loop_1_io_InLiveIn_8_valid),
    .io_InLiveIn_8_bits_predicate(Loop_1_io_InLiveIn_8_bits_predicate),
    .io_InLiveIn_8_bits_taskID(Loop_1_io_InLiveIn_8_bits_taskID),
    .io_InLiveIn_8_bits_data(Loop_1_io_InLiveIn_8_bits_data),
    .io_InLiveIn_9_ready(Loop_1_io_InLiveIn_9_ready),
    .io_InLiveIn_9_valid(Loop_1_io_InLiveIn_9_valid),
    .io_InLiveIn_9_bits_predicate(Loop_1_io_InLiveIn_9_bits_predicate),
    .io_InLiveIn_9_bits_taskID(Loop_1_io_InLiveIn_9_bits_taskID),
    .io_InLiveIn_9_bits_data(Loop_1_io_InLiveIn_9_bits_data),
    .io_InLiveIn_10_ready(Loop_1_io_InLiveIn_10_ready),
    .io_InLiveIn_10_valid(Loop_1_io_InLiveIn_10_valid),
    .io_InLiveIn_10_bits_predicate(Loop_1_io_InLiveIn_10_bits_predicate),
    .io_InLiveIn_10_bits_taskID(Loop_1_io_InLiveIn_10_bits_taskID),
    .io_InLiveIn_10_bits_data(Loop_1_io_InLiveIn_10_bits_data),
    .io_InLiveIn_11_ready(Loop_1_io_InLiveIn_11_ready),
    .io_InLiveIn_11_valid(Loop_1_io_InLiveIn_11_valid),
    .io_InLiveIn_11_bits_predicate(Loop_1_io_InLiveIn_11_bits_predicate),
    .io_InLiveIn_11_bits_taskID(Loop_1_io_InLiveIn_11_bits_taskID),
    .io_InLiveIn_11_bits_data(Loop_1_io_InLiveIn_11_bits_data),
    .io_InLiveIn_12_ready(Loop_1_io_InLiveIn_12_ready),
    .io_InLiveIn_12_valid(Loop_1_io_InLiveIn_12_valid),
    .io_InLiveIn_12_bits_predicate(Loop_1_io_InLiveIn_12_bits_predicate),
    .io_InLiveIn_12_bits_taskID(Loop_1_io_InLiveIn_12_bits_taskID),
    .io_InLiveIn_12_bits_data(Loop_1_io_InLiveIn_12_bits_data),
    .io_OutLiveIn_field12_0_ready(Loop_1_io_OutLiveIn_field12_0_ready),
    .io_OutLiveIn_field12_0_valid(Loop_1_io_OutLiveIn_field12_0_valid),
    .io_OutLiveIn_field12_0_bits_predicate(Loop_1_io_OutLiveIn_field12_0_bits_predicate),
    .io_OutLiveIn_field12_0_bits_taskID(Loop_1_io_OutLiveIn_field12_0_bits_taskID),
    .io_OutLiveIn_field12_0_bits_data(Loop_1_io_OutLiveIn_field12_0_bits_data),
    .io_OutLiveIn_field11_0_ready(Loop_1_io_OutLiveIn_field11_0_ready),
    .io_OutLiveIn_field11_0_valid(Loop_1_io_OutLiveIn_field11_0_valid),
    .io_OutLiveIn_field11_0_bits_predicate(Loop_1_io_OutLiveIn_field11_0_bits_predicate),
    .io_OutLiveIn_field11_0_bits_taskID(Loop_1_io_OutLiveIn_field11_0_bits_taskID),
    .io_OutLiveIn_field11_0_bits_data(Loop_1_io_OutLiveIn_field11_0_bits_data),
    .io_OutLiveIn_field10_0_ready(Loop_1_io_OutLiveIn_field10_0_ready),
    .io_OutLiveIn_field10_0_valid(Loop_1_io_OutLiveIn_field10_0_valid),
    .io_OutLiveIn_field10_0_bits_predicate(Loop_1_io_OutLiveIn_field10_0_bits_predicate),
    .io_OutLiveIn_field10_0_bits_taskID(Loop_1_io_OutLiveIn_field10_0_bits_taskID),
    .io_OutLiveIn_field10_0_bits_data(Loop_1_io_OutLiveIn_field10_0_bits_data),
    .io_OutLiveIn_field9_0_ready(Loop_1_io_OutLiveIn_field9_0_ready),
    .io_OutLiveIn_field9_0_valid(Loop_1_io_OutLiveIn_field9_0_valid),
    .io_OutLiveIn_field9_0_bits_predicate(Loop_1_io_OutLiveIn_field9_0_bits_predicate),
    .io_OutLiveIn_field9_0_bits_taskID(Loop_1_io_OutLiveIn_field9_0_bits_taskID),
    .io_OutLiveIn_field9_0_bits_data(Loop_1_io_OutLiveIn_field9_0_bits_data),
    .io_OutLiveIn_field8_0_ready(Loop_1_io_OutLiveIn_field8_0_ready),
    .io_OutLiveIn_field8_0_valid(Loop_1_io_OutLiveIn_field8_0_valid),
    .io_OutLiveIn_field8_0_bits_predicate(Loop_1_io_OutLiveIn_field8_0_bits_predicate),
    .io_OutLiveIn_field8_0_bits_taskID(Loop_1_io_OutLiveIn_field8_0_bits_taskID),
    .io_OutLiveIn_field8_0_bits_data(Loop_1_io_OutLiveIn_field8_0_bits_data),
    .io_OutLiveIn_field7_0_ready(Loop_1_io_OutLiveIn_field7_0_ready),
    .io_OutLiveIn_field7_0_valid(Loop_1_io_OutLiveIn_field7_0_valid),
    .io_OutLiveIn_field7_0_bits_predicate(Loop_1_io_OutLiveIn_field7_0_bits_predicate),
    .io_OutLiveIn_field7_0_bits_taskID(Loop_1_io_OutLiveIn_field7_0_bits_taskID),
    .io_OutLiveIn_field7_0_bits_data(Loop_1_io_OutLiveIn_field7_0_bits_data),
    .io_OutLiveIn_field6_0_ready(Loop_1_io_OutLiveIn_field6_0_ready),
    .io_OutLiveIn_field6_0_valid(Loop_1_io_OutLiveIn_field6_0_valid),
    .io_OutLiveIn_field6_0_bits_predicate(Loop_1_io_OutLiveIn_field6_0_bits_predicate),
    .io_OutLiveIn_field6_0_bits_taskID(Loop_1_io_OutLiveIn_field6_0_bits_taskID),
    .io_OutLiveIn_field6_0_bits_data(Loop_1_io_OutLiveIn_field6_0_bits_data),
    .io_OutLiveIn_field5_0_ready(Loop_1_io_OutLiveIn_field5_0_ready),
    .io_OutLiveIn_field5_0_valid(Loop_1_io_OutLiveIn_field5_0_valid),
    .io_OutLiveIn_field5_0_bits_predicate(Loop_1_io_OutLiveIn_field5_0_bits_predicate),
    .io_OutLiveIn_field5_0_bits_taskID(Loop_1_io_OutLiveIn_field5_0_bits_taskID),
    .io_OutLiveIn_field5_0_bits_data(Loop_1_io_OutLiveIn_field5_0_bits_data),
    .io_OutLiveIn_field4_0_ready(Loop_1_io_OutLiveIn_field4_0_ready),
    .io_OutLiveIn_field4_0_valid(Loop_1_io_OutLiveIn_field4_0_valid),
    .io_OutLiveIn_field4_0_bits_taskID(Loop_1_io_OutLiveIn_field4_0_bits_taskID),
    .io_OutLiveIn_field4_0_bits_data(Loop_1_io_OutLiveIn_field4_0_bits_data),
    .io_OutLiveIn_field3_0_ready(Loop_1_io_OutLiveIn_field3_0_ready),
    .io_OutLiveIn_field3_0_valid(Loop_1_io_OutLiveIn_field3_0_valid),
    .io_OutLiveIn_field3_0_bits_predicate(Loop_1_io_OutLiveIn_field3_0_bits_predicate),
    .io_OutLiveIn_field3_0_bits_taskID(Loop_1_io_OutLiveIn_field3_0_bits_taskID),
    .io_OutLiveIn_field3_0_bits_data(Loop_1_io_OutLiveIn_field3_0_bits_data),
    .io_OutLiveIn_field2_0_ready(Loop_1_io_OutLiveIn_field2_0_ready),
    .io_OutLiveIn_field2_0_valid(Loop_1_io_OutLiveIn_field2_0_valid),
    .io_OutLiveIn_field2_0_bits_taskID(Loop_1_io_OutLiveIn_field2_0_bits_taskID),
    .io_OutLiveIn_field2_0_bits_data(Loop_1_io_OutLiveIn_field2_0_bits_data),
    .io_OutLiveIn_field1_0_ready(Loop_1_io_OutLiveIn_field1_0_ready),
    .io_OutLiveIn_field1_0_valid(Loop_1_io_OutLiveIn_field1_0_valid),
    .io_OutLiveIn_field1_0_bits_data(Loop_1_io_OutLiveIn_field1_0_bits_data),
    .io_OutLiveIn_field1_1_ready(Loop_1_io_OutLiveIn_field1_1_ready),
    .io_OutLiveIn_field1_1_valid(Loop_1_io_OutLiveIn_field1_1_valid),
    .io_OutLiveIn_field1_1_bits_data(Loop_1_io_OutLiveIn_field1_1_bits_data),
    .io_OutLiveIn_field1_2_ready(Loop_1_io_OutLiveIn_field1_2_ready),
    .io_OutLiveIn_field1_2_valid(Loop_1_io_OutLiveIn_field1_2_valid),
    .io_OutLiveIn_field1_2_bits_data(Loop_1_io_OutLiveIn_field1_2_bits_data),
    .io_OutLiveIn_field0_0_ready(Loop_1_io_OutLiveIn_field0_0_ready),
    .io_OutLiveIn_field0_0_valid(Loop_1_io_OutLiveIn_field0_0_valid),
    .io_OutLiveIn_field0_0_bits_data(Loop_1_io_OutLiveIn_field0_0_bits_data),
    .io_OutLiveIn_field0_1_ready(Loop_1_io_OutLiveIn_field0_1_ready),
    .io_OutLiveIn_field0_1_valid(Loop_1_io_OutLiveIn_field0_1_valid),
    .io_OutLiveIn_field0_1_bits_data(Loop_1_io_OutLiveIn_field0_1_bits_data),
    .io_OutLiveIn_field0_2_ready(Loop_1_io_OutLiveIn_field0_2_ready),
    .io_OutLiveIn_field0_2_valid(Loop_1_io_OutLiveIn_field0_2_valid),
    .io_OutLiveIn_field0_2_bits_data(Loop_1_io_OutLiveIn_field0_2_bits_data),
    .io_activate_loop_start_ready(Loop_1_io_activate_loop_start_ready),
    .io_activate_loop_start_valid(Loop_1_io_activate_loop_start_valid),
    .io_activate_loop_start_bits_taskID(Loop_1_io_activate_loop_start_bits_taskID),
    .io_activate_loop_start_bits_control(Loop_1_io_activate_loop_start_bits_control),
    .io_activate_loop_back_ready(Loop_1_io_activate_loop_back_ready),
    .io_activate_loop_back_valid(Loop_1_io_activate_loop_back_valid),
    .io_activate_loop_back_bits_taskID(Loop_1_io_activate_loop_back_bits_taskID),
    .io_activate_loop_back_bits_control(Loop_1_io_activate_loop_back_bits_control),
    .io_loopBack_0_ready(Loop_1_io_loopBack_0_ready),
    .io_loopBack_0_valid(Loop_1_io_loopBack_0_valid),
    .io_loopBack_0_bits_taskID(Loop_1_io_loopBack_0_bits_taskID),
    .io_loopBack_0_bits_control(Loop_1_io_loopBack_0_bits_control),
    .io_loopFinish_0_ready(Loop_1_io_loopFinish_0_ready),
    .io_loopFinish_0_valid(Loop_1_io_loopFinish_0_valid),
    .io_loopFinish_0_bits_control(Loop_1_io_loopFinish_0_bits_control),
    .io_CarryDepenIn_0_ready(Loop_1_io_CarryDepenIn_0_ready),
    .io_CarryDepenIn_0_valid(Loop_1_io_CarryDepenIn_0_valid),
    .io_CarryDepenIn_0_bits_taskID(Loop_1_io_CarryDepenIn_0_bits_taskID),
    .io_CarryDepenIn_0_bits_data(Loop_1_io_CarryDepenIn_0_bits_data),
    .io_CarryDepenOut_field0_0_ready(Loop_1_io_CarryDepenOut_field0_0_ready),
    .io_CarryDepenOut_field0_0_valid(Loop_1_io_CarryDepenOut_field0_0_valid),
    .io_CarryDepenOut_field0_0_bits_taskID(Loop_1_io_CarryDepenOut_field0_0_bits_taskID),
    .io_CarryDepenOut_field0_0_bits_data(Loop_1_io_CarryDepenOut_field0_0_bits_data),
    .io_loopExit_0_ready(Loop_1_io_loopExit_0_ready),
    .io_loopExit_0_valid(Loop_1_io_loopExit_0_valid),
    .io_loopExit_0_bits_taskID(Loop_1_io_loopExit_0_bits_taskID),
    .io_loopExit_0_bits_control(Loop_1_io_loopExit_0_bits_control)
  );
  BasicBlockNoMaskFastNode bb_entry0 ( // @[extracted_function_conv.scala 72:25]
    .clock(bb_entry0_clock),
    .reset(bb_entry0_reset),
    .io_predicateIn_0_ready(bb_entry0_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_entry0_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_entry0_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_entry0_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_entry0_io_Out_0_ready),
    .io_Out_0_valid(bb_entry0_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_entry0_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_entry0_io_Out_1_ready),
    .io_Out_1_valid(bb_entry0_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_entry0_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_entry0_io_Out_2_ready),
    .io_Out_2_valid(bb_entry0_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_entry0_io_Out_2_bits_taskID),
    .io_Out_3_ready(bb_entry0_io_Out_3_ready),
    .io_Out_3_valid(bb_entry0_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_entry0_io_Out_3_bits_taskID),
    .io_Out_4_ready(bb_entry0_io_Out_4_ready),
    .io_Out_4_valid(bb_entry0_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_entry0_io_Out_4_bits_taskID),
    .io_Out_5_ready(bb_entry0_io_Out_5_ready),
    .io_Out_5_valid(bb_entry0_io_Out_5_valid),
    .io_Out_5_bits_taskID(bb_entry0_io_Out_5_bits_taskID),
    .io_Out_6_ready(bb_entry0_io_Out_6_ready),
    .io_Out_6_valid(bb_entry0_io_Out_6_valid),
    .io_Out_6_bits_taskID(bb_entry0_io_Out_6_bits_taskID),
    .io_Out_7_ready(bb_entry0_io_Out_7_ready),
    .io_Out_7_valid(bb_entry0_io_Out_7_valid),
    .io_Out_7_bits_taskID(bb_entry0_io_Out_7_bits_taskID),
    .io_Out_8_ready(bb_entry0_io_Out_8_ready),
    .io_Out_8_valid(bb_entry0_io_Out_8_valid),
    .io_Out_8_bits_taskID(bb_entry0_io_Out_8_bits_taskID),
    .io_Out_8_bits_control(bb_entry0_io_Out_8_bits_control),
    .io_Out_9_ready(bb_entry0_io_Out_9_ready),
    .io_Out_9_valid(bb_entry0_io_Out_9_valid),
    .io_Out_9_bits_taskID(bb_entry0_io_Out_9_bits_taskID),
    .io_Out_9_bits_control(bb_entry0_io_Out_9_bits_control),
    .io_Out_10_ready(bb_entry0_io_Out_10_ready),
    .io_Out_10_valid(bb_entry0_io_Out_10_valid),
    .io_Out_10_bits_taskID(bb_entry0_io_Out_10_bits_taskID),
    .io_Out_10_bits_control(bb_entry0_io_Out_10_bits_control),
    .io_Out_11_ready(bb_entry0_io_Out_11_ready),
    .io_Out_11_valid(bb_entry0_io_Out_11_valid),
    .io_Out_11_bits_taskID(bb_entry0_io_Out_11_bits_taskID),
    .io_Out_11_bits_control(bb_entry0_io_Out_11_bits_control),
    .io_Out_12_ready(bb_entry0_io_Out_12_ready),
    .io_Out_12_valid(bb_entry0_io_Out_12_valid),
    .io_Out_12_bits_taskID(bb_entry0_io_Out_12_bits_taskID),
    .io_Out_12_bits_control(bb_entry0_io_Out_12_bits_control),
    .io_Out_13_ready(bb_entry0_io_Out_13_ready),
    .io_Out_13_valid(bb_entry0_io_Out_13_valid),
    .io_Out_13_bits_taskID(bb_entry0_io_Out_13_bits_taskID),
    .io_Out_13_bits_control(bb_entry0_io_Out_13_bits_control),
    .io_Out_14_ready(bb_entry0_io_Out_14_ready),
    .io_Out_14_valid(bb_entry0_io_Out_14_valid),
    .io_Out_14_bits_taskID(bb_entry0_io_Out_14_bits_taskID),
    .io_Out_14_bits_control(bb_entry0_io_Out_14_bits_control),
    .io_Out_15_ready(bb_entry0_io_Out_15_ready),
    .io_Out_15_valid(bb_entry0_io_Out_15_valid),
    .io_Out_15_bits_taskID(bb_entry0_io_Out_15_bits_taskID),
    .io_Out_15_bits_control(bb_entry0_io_Out_15_bits_control),
    .io_Out_16_ready(bb_entry0_io_Out_16_ready),
    .io_Out_16_valid(bb_entry0_io_Out_16_valid),
    .io_Out_16_bits_taskID(bb_entry0_io_Out_16_bits_taskID),
    .io_Out_16_bits_control(bb_entry0_io_Out_16_bits_control),
    .io_Out_17_ready(bb_entry0_io_Out_17_ready),
    .io_Out_17_valid(bb_entry0_io_Out_17_valid),
    .io_Out_17_bits_taskID(bb_entry0_io_Out_17_bits_taskID),
    .io_Out_17_bits_control(bb_entry0_io_Out_17_bits_control),
    .io_Out_18_ready(bb_entry0_io_Out_18_ready),
    .io_Out_18_valid(bb_entry0_io_Out_18_valid),
    .io_Out_18_bits_taskID(bb_entry0_io_Out_18_bits_taskID),
    .io_Out_18_bits_control(bb_entry0_io_Out_18_bits_control)
  );
  BasicBlockNoMaskFastNode_1 bb_for_cond_cleanup1 ( // @[extracted_function_conv.scala 74:36]
    .clock(bb_for_cond_cleanup1_clock),
    .reset(bb_for_cond_cleanup1_reset),
    .io_predicateIn_0_ready(bb_for_cond_cleanup1_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup1_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup1_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup1_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_cond_cleanup1_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup1_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup1_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(bb_for_cond_cleanup1_io_Out_0_bits_control)
  );
  BasicBlockNode bb_for_body2 ( // @[extracted_function_conv.scala 76:28]
    .clock(bb_for_body2_clock),
    .reset(bb_for_body2_reset),
    .io_MaskBB_0_ready(bb_for_body2_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body2_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body2_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_for_body2_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body2_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body2_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_body2_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body2_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body2_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_for_body2_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body2_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body2_io_Out_2_bits_taskID),
    .io_Out_3_ready(bb_for_body2_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body2_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_body2_io_Out_3_bits_taskID),
    .io_Out_4_ready(bb_for_body2_io_Out_4_ready),
    .io_Out_4_valid(bb_for_body2_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_body2_io_Out_4_bits_taskID),
    .io_Out_5_ready(bb_for_body2_io_Out_5_ready),
    .io_Out_5_valid(bb_for_body2_io_Out_5_valid),
    .io_Out_5_bits_control(bb_for_body2_io_Out_5_bits_control),
    .io_Out_6_ready(bb_for_body2_io_Out_6_ready),
    .io_Out_6_valid(bb_for_body2_io_Out_6_valid),
    .io_Out_6_bits_taskID(bb_for_body2_io_Out_6_bits_taskID),
    .io_Out_6_bits_control(bb_for_body2_io_Out_6_bits_control),
    .io_Out_7_ready(bb_for_body2_io_Out_7_ready),
    .io_Out_7_valid(bb_for_body2_io_Out_7_valid),
    .io_Out_7_bits_taskID(bb_for_body2_io_Out_7_bits_taskID),
    .io_Out_7_bits_control(bb_for_body2_io_Out_7_bits_control),
    .io_Out_8_ready(bb_for_body2_io_Out_8_ready),
    .io_Out_8_valid(bb_for_body2_io_Out_8_valid),
    .io_Out_8_bits_taskID(bb_for_body2_io_Out_8_bits_taskID),
    .io_Out_8_bits_control(bb_for_body2_io_Out_8_bits_control),
    .io_Out_9_ready(bb_for_body2_io_Out_9_ready),
    .io_Out_9_valid(bb_for_body2_io_Out_9_valid),
    .io_Out_9_bits_taskID(bb_for_body2_io_Out_9_bits_taskID),
    .io_Out_9_bits_control(bb_for_body2_io_Out_9_bits_control),
    .io_Out_10_ready(bb_for_body2_io_Out_10_ready),
    .io_Out_10_valid(bb_for_body2_io_Out_10_valid),
    .io_Out_10_bits_taskID(bb_for_body2_io_Out_10_bits_taskID),
    .io_Out_10_bits_control(bb_for_body2_io_Out_10_bits_control),
    .io_Out_11_ready(bb_for_body2_io_Out_11_ready),
    .io_Out_11_valid(bb_for_body2_io_Out_11_valid),
    .io_Out_11_bits_taskID(bb_for_body2_io_Out_11_bits_taskID),
    .io_Out_11_bits_control(bb_for_body2_io_Out_11_bits_control),
    .io_Out_12_ready(bb_for_body2_io_Out_12_ready),
    .io_Out_12_valid(bb_for_body2_io_Out_12_valid),
    .io_Out_12_bits_taskID(bb_for_body2_io_Out_12_bits_taskID),
    .io_Out_12_bits_control(bb_for_body2_io_Out_12_bits_control),
    .io_Out_13_ready(bb_for_body2_io_Out_13_ready),
    .io_Out_13_valid(bb_for_body2_io_Out_13_valid),
    .io_Out_13_bits_taskID(bb_for_body2_io_Out_13_bits_taskID),
    .io_Out_13_bits_control(bb_for_body2_io_Out_13_bits_control),
    .io_Out_14_ready(bb_for_body2_io_Out_14_ready),
    .io_Out_14_valid(bb_for_body2_io_Out_14_valid),
    .io_Out_14_bits_taskID(bb_for_body2_io_Out_14_bits_taskID),
    .io_Out_14_bits_control(bb_for_body2_io_Out_14_bits_control),
    .io_Out_15_ready(bb_for_body2_io_Out_15_ready),
    .io_Out_15_valid(bb_for_body2_io_Out_15_valid),
    .io_Out_15_bits_taskID(bb_for_body2_io_Out_15_bits_taskID),
    .io_Out_15_bits_control(bb_for_body2_io_Out_15_bits_control),
    .io_predicateIn_0_ready(bb_for_body2_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body2_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body2_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body2_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body2_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body2_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body2_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body2_io_predicateIn_1_bits_control)
  );
  BasicBlockNoMaskFastNode_2 bb_for_cond_cleanup113 ( // @[extracted_function_conv.scala 78:38]
    .clock(bb_for_cond_cleanup113_clock),
    .reset(bb_for_cond_cleanup113_reset),
    .io_predicateIn_0_ready(bb_for_cond_cleanup113_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_cond_cleanup113_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_cond_cleanup113_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_cond_cleanup113_io_predicateIn_0_bits_control),
    .io_Out_0_ready(bb_for_cond_cleanup113_io_Out_0_ready),
    .io_Out_0_valid(bb_for_cond_cleanup113_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_cond_cleanup113_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_cond_cleanup113_io_Out_1_ready),
    .io_Out_1_valid(bb_for_cond_cleanup113_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_cond_cleanup113_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_for_cond_cleanup113_io_Out_2_ready),
    .io_Out_2_valid(bb_for_cond_cleanup113_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_cond_cleanup113_io_Out_2_bits_taskID),
    .io_Out_2_bits_control(bb_for_cond_cleanup113_io_Out_2_bits_control),
    .io_Out_3_ready(bb_for_cond_cleanup113_io_Out_3_ready),
    .io_Out_3_valid(bb_for_cond_cleanup113_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_cond_cleanup113_io_Out_3_bits_taskID),
    .io_Out_3_bits_control(bb_for_cond_cleanup113_io_Out_3_bits_control),
    .io_Out_4_ready(bb_for_cond_cleanup113_io_Out_4_ready),
    .io_Out_4_valid(bb_for_cond_cleanup113_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_cond_cleanup113_io_Out_4_bits_taskID),
    .io_Out_4_bits_control(bb_for_cond_cleanup113_io_Out_4_bits_control)
  );
  BasicBlockNode_1 bb_for_body124 ( // @[extracted_function_conv.scala 80:30]
    .clock(bb_for_body124_clock),
    .reset(bb_for_body124_reset),
    .io_MaskBB_0_ready(bb_for_body124_io_MaskBB_0_ready),
    .io_MaskBB_0_valid(bb_for_body124_io_MaskBB_0_valid),
    .io_MaskBB_0_bits(bb_for_body124_io_MaskBB_0_bits),
    .io_Out_0_ready(bb_for_body124_io_Out_0_ready),
    .io_Out_0_valid(bb_for_body124_io_Out_0_valid),
    .io_Out_0_bits_taskID(bb_for_body124_io_Out_0_bits_taskID),
    .io_Out_1_ready(bb_for_body124_io_Out_1_ready),
    .io_Out_1_valid(bb_for_body124_io_Out_1_valid),
    .io_Out_1_bits_taskID(bb_for_body124_io_Out_1_bits_taskID),
    .io_Out_2_ready(bb_for_body124_io_Out_2_ready),
    .io_Out_2_valid(bb_for_body124_io_Out_2_valid),
    .io_Out_2_bits_taskID(bb_for_body124_io_Out_2_bits_taskID),
    .io_Out_3_ready(bb_for_body124_io_Out_3_ready),
    .io_Out_3_valid(bb_for_body124_io_Out_3_valid),
    .io_Out_3_bits_taskID(bb_for_body124_io_Out_3_bits_taskID),
    .io_Out_4_ready(bb_for_body124_io_Out_4_ready),
    .io_Out_4_valid(bb_for_body124_io_Out_4_valid),
    .io_Out_4_bits_taskID(bb_for_body124_io_Out_4_bits_taskID),
    .io_Out_5_ready(bb_for_body124_io_Out_5_ready),
    .io_Out_5_valid(bb_for_body124_io_Out_5_valid),
    .io_Out_5_bits_taskID(bb_for_body124_io_Out_5_bits_taskID),
    .io_Out_6_ready(bb_for_body124_io_Out_6_ready),
    .io_Out_6_valid(bb_for_body124_io_Out_6_valid),
    .io_Out_6_bits_taskID(bb_for_body124_io_Out_6_bits_taskID),
    .io_Out_7_ready(bb_for_body124_io_Out_7_ready),
    .io_Out_7_valid(bb_for_body124_io_Out_7_valid),
    .io_Out_7_bits_taskID(bb_for_body124_io_Out_7_bits_taskID),
    .io_Out_8_ready(bb_for_body124_io_Out_8_ready),
    .io_Out_8_valid(bb_for_body124_io_Out_8_valid),
    .io_Out_8_bits_taskID(bb_for_body124_io_Out_8_bits_taskID),
    .io_Out_9_ready(bb_for_body124_io_Out_9_ready),
    .io_Out_9_valid(bb_for_body124_io_Out_9_valid),
    .io_Out_9_bits_taskID(bb_for_body124_io_Out_9_bits_taskID),
    .io_Out_10_ready(bb_for_body124_io_Out_10_ready),
    .io_Out_10_valid(bb_for_body124_io_Out_10_valid),
    .io_Out_10_bits_taskID(bb_for_body124_io_Out_10_bits_taskID),
    .io_Out_11_ready(bb_for_body124_io_Out_11_ready),
    .io_Out_11_valid(bb_for_body124_io_Out_11_valid),
    .io_Out_11_bits_control(bb_for_body124_io_Out_11_bits_control),
    .io_Out_12_ready(bb_for_body124_io_Out_12_ready),
    .io_Out_12_valid(bb_for_body124_io_Out_12_valid),
    .io_Out_12_bits_taskID(bb_for_body124_io_Out_12_bits_taskID),
    .io_Out_12_bits_control(bb_for_body124_io_Out_12_bits_control),
    .io_Out_13_ready(bb_for_body124_io_Out_13_ready),
    .io_Out_13_valid(bb_for_body124_io_Out_13_valid),
    .io_Out_13_bits_taskID(bb_for_body124_io_Out_13_bits_taskID),
    .io_Out_13_bits_control(bb_for_body124_io_Out_13_bits_control),
    .io_Out_14_ready(bb_for_body124_io_Out_14_ready),
    .io_Out_14_valid(bb_for_body124_io_Out_14_valid),
    .io_Out_14_bits_taskID(bb_for_body124_io_Out_14_bits_taskID),
    .io_Out_14_bits_control(bb_for_body124_io_Out_14_bits_control),
    .io_Out_15_ready(bb_for_body124_io_Out_15_ready),
    .io_Out_15_valid(bb_for_body124_io_Out_15_valid),
    .io_Out_15_bits_taskID(bb_for_body124_io_Out_15_bits_taskID),
    .io_Out_15_bits_control(bb_for_body124_io_Out_15_bits_control),
    .io_Out_16_ready(bb_for_body124_io_Out_16_ready),
    .io_Out_16_valid(bb_for_body124_io_Out_16_valid),
    .io_Out_16_bits_taskID(bb_for_body124_io_Out_16_bits_taskID),
    .io_Out_16_bits_control(bb_for_body124_io_Out_16_bits_control),
    .io_Out_17_ready(bb_for_body124_io_Out_17_ready),
    .io_Out_17_valid(bb_for_body124_io_Out_17_valid),
    .io_Out_17_bits_taskID(bb_for_body124_io_Out_17_bits_taskID),
    .io_Out_17_bits_control(bb_for_body124_io_Out_17_bits_control),
    .io_Out_18_ready(bb_for_body124_io_Out_18_ready),
    .io_Out_18_valid(bb_for_body124_io_Out_18_valid),
    .io_Out_18_bits_taskID(bb_for_body124_io_Out_18_bits_taskID),
    .io_Out_18_bits_control(bb_for_body124_io_Out_18_bits_control),
    .io_Out_19_ready(bb_for_body124_io_Out_19_ready),
    .io_Out_19_valid(bb_for_body124_io_Out_19_valid),
    .io_Out_19_bits_taskID(bb_for_body124_io_Out_19_bits_taskID),
    .io_Out_19_bits_control(bb_for_body124_io_Out_19_bits_control),
    .io_Out_20_ready(bb_for_body124_io_Out_20_ready),
    .io_Out_20_valid(bb_for_body124_io_Out_20_valid),
    .io_Out_20_bits_taskID(bb_for_body124_io_Out_20_bits_taskID),
    .io_Out_20_bits_control(bb_for_body124_io_Out_20_bits_control),
    .io_Out_21_ready(bb_for_body124_io_Out_21_ready),
    .io_Out_21_valid(bb_for_body124_io_Out_21_valid),
    .io_Out_21_bits_taskID(bb_for_body124_io_Out_21_bits_taskID),
    .io_Out_22_ready(bb_for_body124_io_Out_22_ready),
    .io_Out_22_valid(bb_for_body124_io_Out_22_valid),
    .io_Out_22_bits_taskID(bb_for_body124_io_Out_22_bits_taskID),
    .io_Out_22_bits_control(bb_for_body124_io_Out_22_bits_control),
    .io_Out_23_ready(bb_for_body124_io_Out_23_ready),
    .io_Out_23_valid(bb_for_body124_io_Out_23_valid),
    .io_Out_23_bits_taskID(bb_for_body124_io_Out_23_bits_taskID),
    .io_Out_23_bits_control(bb_for_body124_io_Out_23_bits_control),
    .io_Out_24_ready(bb_for_body124_io_Out_24_ready),
    .io_Out_24_valid(bb_for_body124_io_Out_24_valid),
    .io_Out_24_bits_taskID(bb_for_body124_io_Out_24_bits_taskID),
    .io_Out_24_bits_control(bb_for_body124_io_Out_24_bits_control),
    .io_Out_25_ready(bb_for_body124_io_Out_25_ready),
    .io_Out_25_valid(bb_for_body124_io_Out_25_valid),
    .io_Out_25_bits_taskID(bb_for_body124_io_Out_25_bits_taskID),
    .io_Out_25_bits_control(bb_for_body124_io_Out_25_bits_control),
    .io_Out_26_ready(bb_for_body124_io_Out_26_ready),
    .io_Out_26_valid(bb_for_body124_io_Out_26_valid),
    .io_Out_26_bits_taskID(bb_for_body124_io_Out_26_bits_taskID),
    .io_Out_26_bits_control(bb_for_body124_io_Out_26_bits_control),
    .io_Out_27_ready(bb_for_body124_io_Out_27_ready),
    .io_Out_27_valid(bb_for_body124_io_Out_27_valid),
    .io_Out_27_bits_taskID(bb_for_body124_io_Out_27_bits_taskID),
    .io_Out_27_bits_control(bb_for_body124_io_Out_27_bits_control),
    .io_Out_28_ready(bb_for_body124_io_Out_28_ready),
    .io_Out_28_valid(bb_for_body124_io_Out_28_valid),
    .io_Out_28_bits_taskID(bb_for_body124_io_Out_28_bits_taskID),
    .io_Out_28_bits_control(bb_for_body124_io_Out_28_bits_control),
    .io_Out_29_ready(bb_for_body124_io_Out_29_ready),
    .io_Out_29_valid(bb_for_body124_io_Out_29_valid),
    .io_Out_29_bits_taskID(bb_for_body124_io_Out_29_bits_taskID),
    .io_Out_30_ready(bb_for_body124_io_Out_30_ready),
    .io_Out_30_valid(bb_for_body124_io_Out_30_valid),
    .io_Out_30_bits_taskID(bb_for_body124_io_Out_30_bits_taskID),
    .io_Out_30_bits_control(bb_for_body124_io_Out_30_bits_control),
    .io_Out_31_ready(bb_for_body124_io_Out_31_ready),
    .io_Out_31_valid(bb_for_body124_io_Out_31_valid),
    .io_Out_31_bits_taskID(bb_for_body124_io_Out_31_bits_taskID),
    .io_Out_31_bits_control(bb_for_body124_io_Out_31_bits_control),
    .io_Out_32_ready(bb_for_body124_io_Out_32_ready),
    .io_Out_32_valid(bb_for_body124_io_Out_32_valid),
    .io_Out_32_bits_taskID(bb_for_body124_io_Out_32_bits_taskID),
    .io_Out_32_bits_control(bb_for_body124_io_Out_32_bits_control),
    .io_Out_33_ready(bb_for_body124_io_Out_33_ready),
    .io_Out_33_valid(bb_for_body124_io_Out_33_valid),
    .io_Out_33_bits_taskID(bb_for_body124_io_Out_33_bits_taskID),
    .io_Out_33_bits_control(bb_for_body124_io_Out_33_bits_control),
    .io_Out_34_ready(bb_for_body124_io_Out_34_ready),
    .io_Out_34_valid(bb_for_body124_io_Out_34_valid),
    .io_Out_34_bits_taskID(bb_for_body124_io_Out_34_bits_taskID),
    .io_Out_34_bits_control(bb_for_body124_io_Out_34_bits_control),
    .io_Out_35_ready(bb_for_body124_io_Out_35_ready),
    .io_Out_35_valid(bb_for_body124_io_Out_35_valid),
    .io_Out_35_bits_taskID(bb_for_body124_io_Out_35_bits_taskID),
    .io_Out_35_bits_control(bb_for_body124_io_Out_35_bits_control),
    .io_Out_36_ready(bb_for_body124_io_Out_36_ready),
    .io_Out_36_valid(bb_for_body124_io_Out_36_valid),
    .io_Out_36_bits_taskID(bb_for_body124_io_Out_36_bits_taskID),
    .io_Out_36_bits_control(bb_for_body124_io_Out_36_bits_control),
    .io_Out_37_ready(bb_for_body124_io_Out_37_ready),
    .io_Out_37_valid(bb_for_body124_io_Out_37_valid),
    .io_Out_37_bits_taskID(bb_for_body124_io_Out_37_bits_taskID),
    .io_Out_38_ready(bb_for_body124_io_Out_38_ready),
    .io_Out_38_valid(bb_for_body124_io_Out_38_valid),
    .io_Out_38_bits_taskID(bb_for_body124_io_Out_38_bits_taskID),
    .io_Out_38_bits_control(bb_for_body124_io_Out_38_bits_control),
    .io_Out_39_ready(bb_for_body124_io_Out_39_ready),
    .io_Out_39_valid(bb_for_body124_io_Out_39_valid),
    .io_Out_39_bits_taskID(bb_for_body124_io_Out_39_bits_taskID),
    .io_Out_39_bits_control(bb_for_body124_io_Out_39_bits_control),
    .io_Out_40_ready(bb_for_body124_io_Out_40_ready),
    .io_Out_40_valid(bb_for_body124_io_Out_40_valid),
    .io_Out_40_bits_taskID(bb_for_body124_io_Out_40_bits_taskID),
    .io_Out_40_bits_control(bb_for_body124_io_Out_40_bits_control),
    .io_Out_41_ready(bb_for_body124_io_Out_41_ready),
    .io_Out_41_valid(bb_for_body124_io_Out_41_valid),
    .io_Out_41_bits_taskID(bb_for_body124_io_Out_41_bits_taskID),
    .io_Out_41_bits_control(bb_for_body124_io_Out_41_bits_control),
    .io_Out_42_ready(bb_for_body124_io_Out_42_ready),
    .io_Out_42_valid(bb_for_body124_io_Out_42_valid),
    .io_Out_42_bits_taskID(bb_for_body124_io_Out_42_bits_taskID),
    .io_Out_42_bits_control(bb_for_body124_io_Out_42_bits_control),
    .io_Out_43_ready(bb_for_body124_io_Out_43_ready),
    .io_Out_43_valid(bb_for_body124_io_Out_43_valid),
    .io_Out_43_bits_taskID(bb_for_body124_io_Out_43_bits_taskID),
    .io_Out_43_bits_control(bb_for_body124_io_Out_43_bits_control),
    .io_Out_44_ready(bb_for_body124_io_Out_44_ready),
    .io_Out_44_valid(bb_for_body124_io_Out_44_valid),
    .io_Out_44_bits_taskID(bb_for_body124_io_Out_44_bits_taskID),
    .io_Out_44_bits_control(bb_for_body124_io_Out_44_bits_control),
    .io_Out_45_ready(bb_for_body124_io_Out_45_ready),
    .io_Out_45_valid(bb_for_body124_io_Out_45_valid),
    .io_Out_45_bits_taskID(bb_for_body124_io_Out_45_bits_taskID),
    .io_Out_45_bits_control(bb_for_body124_io_Out_45_bits_control),
    .io_Out_46_ready(bb_for_body124_io_Out_46_ready),
    .io_Out_46_valid(bb_for_body124_io_Out_46_valid),
    .io_Out_46_bits_taskID(bb_for_body124_io_Out_46_bits_taskID),
    .io_Out_47_ready(bb_for_body124_io_Out_47_ready),
    .io_Out_47_valid(bb_for_body124_io_Out_47_valid),
    .io_Out_47_bits_taskID(bb_for_body124_io_Out_47_bits_taskID),
    .io_Out_47_bits_control(bb_for_body124_io_Out_47_bits_control),
    .io_Out_48_ready(bb_for_body124_io_Out_48_ready),
    .io_Out_48_valid(bb_for_body124_io_Out_48_valid),
    .io_Out_48_bits_taskID(bb_for_body124_io_Out_48_bits_taskID),
    .io_Out_48_bits_control(bb_for_body124_io_Out_48_bits_control),
    .io_Out_49_ready(bb_for_body124_io_Out_49_ready),
    .io_Out_49_valid(bb_for_body124_io_Out_49_valid),
    .io_Out_49_bits_taskID(bb_for_body124_io_Out_49_bits_taskID),
    .io_Out_49_bits_control(bb_for_body124_io_Out_49_bits_control),
    .io_Out_50_ready(bb_for_body124_io_Out_50_ready),
    .io_Out_50_valid(bb_for_body124_io_Out_50_valid),
    .io_Out_50_bits_taskID(bb_for_body124_io_Out_50_bits_taskID),
    .io_Out_50_bits_control(bb_for_body124_io_Out_50_bits_control),
    .io_Out_51_ready(bb_for_body124_io_Out_51_ready),
    .io_Out_51_valid(bb_for_body124_io_Out_51_valid),
    .io_Out_51_bits_taskID(bb_for_body124_io_Out_51_bits_taskID),
    .io_Out_51_bits_control(bb_for_body124_io_Out_51_bits_control),
    .io_Out_52_ready(bb_for_body124_io_Out_52_ready),
    .io_Out_52_valid(bb_for_body124_io_Out_52_valid),
    .io_Out_52_bits_taskID(bb_for_body124_io_Out_52_bits_taskID),
    .io_Out_52_bits_control(bb_for_body124_io_Out_52_bits_control),
    .io_Out_53_ready(bb_for_body124_io_Out_53_ready),
    .io_Out_53_valid(bb_for_body124_io_Out_53_valid),
    .io_Out_53_bits_taskID(bb_for_body124_io_Out_53_bits_taskID),
    .io_Out_53_bits_control(bb_for_body124_io_Out_53_bits_control),
    .io_Out_54_ready(bb_for_body124_io_Out_54_ready),
    .io_Out_54_valid(bb_for_body124_io_Out_54_valid),
    .io_Out_54_bits_taskID(bb_for_body124_io_Out_54_bits_taskID),
    .io_Out_55_ready(bb_for_body124_io_Out_55_ready),
    .io_Out_55_valid(bb_for_body124_io_Out_55_valid),
    .io_Out_55_bits_taskID(bb_for_body124_io_Out_55_bits_taskID),
    .io_Out_55_bits_control(bb_for_body124_io_Out_55_bits_control),
    .io_Out_56_ready(bb_for_body124_io_Out_56_ready),
    .io_Out_56_valid(bb_for_body124_io_Out_56_valid),
    .io_Out_56_bits_taskID(bb_for_body124_io_Out_56_bits_taskID),
    .io_Out_56_bits_control(bb_for_body124_io_Out_56_bits_control),
    .io_Out_57_ready(bb_for_body124_io_Out_57_ready),
    .io_Out_57_valid(bb_for_body124_io_Out_57_valid),
    .io_Out_57_bits_taskID(bb_for_body124_io_Out_57_bits_taskID),
    .io_Out_57_bits_control(bb_for_body124_io_Out_57_bits_control),
    .io_Out_58_ready(bb_for_body124_io_Out_58_ready),
    .io_Out_58_valid(bb_for_body124_io_Out_58_valid),
    .io_Out_58_bits_taskID(bb_for_body124_io_Out_58_bits_taskID),
    .io_Out_58_bits_control(bb_for_body124_io_Out_58_bits_control),
    .io_Out_59_ready(bb_for_body124_io_Out_59_ready),
    .io_Out_59_valid(bb_for_body124_io_Out_59_valid),
    .io_Out_59_bits_taskID(bb_for_body124_io_Out_59_bits_taskID),
    .io_Out_59_bits_control(bb_for_body124_io_Out_59_bits_control),
    .io_Out_60_ready(bb_for_body124_io_Out_60_ready),
    .io_Out_60_valid(bb_for_body124_io_Out_60_valid),
    .io_Out_60_bits_taskID(bb_for_body124_io_Out_60_bits_taskID),
    .io_Out_60_bits_control(bb_for_body124_io_Out_60_bits_control),
    .io_Out_61_ready(bb_for_body124_io_Out_61_ready),
    .io_Out_61_valid(bb_for_body124_io_Out_61_valid),
    .io_Out_61_bits_taskID(bb_for_body124_io_Out_61_bits_taskID),
    .io_Out_61_bits_control(bb_for_body124_io_Out_61_bits_control),
    .io_Out_62_ready(bb_for_body124_io_Out_62_ready),
    .io_Out_62_valid(bb_for_body124_io_Out_62_valid),
    .io_Out_62_bits_taskID(bb_for_body124_io_Out_62_bits_taskID),
    .io_Out_63_ready(bb_for_body124_io_Out_63_ready),
    .io_Out_63_valid(bb_for_body124_io_Out_63_valid),
    .io_Out_63_bits_taskID(bb_for_body124_io_Out_63_bits_taskID),
    .io_Out_63_bits_control(bb_for_body124_io_Out_63_bits_control),
    .io_Out_64_ready(bb_for_body124_io_Out_64_ready),
    .io_Out_64_valid(bb_for_body124_io_Out_64_valid),
    .io_Out_64_bits_taskID(bb_for_body124_io_Out_64_bits_taskID),
    .io_Out_64_bits_control(bb_for_body124_io_Out_64_bits_control),
    .io_Out_65_ready(bb_for_body124_io_Out_65_ready),
    .io_Out_65_valid(bb_for_body124_io_Out_65_valid),
    .io_Out_65_bits_taskID(bb_for_body124_io_Out_65_bits_taskID),
    .io_Out_65_bits_control(bb_for_body124_io_Out_65_bits_control),
    .io_Out_66_ready(bb_for_body124_io_Out_66_ready),
    .io_Out_66_valid(bb_for_body124_io_Out_66_valid),
    .io_Out_66_bits_taskID(bb_for_body124_io_Out_66_bits_taskID),
    .io_Out_66_bits_control(bb_for_body124_io_Out_66_bits_control),
    .io_Out_67_ready(bb_for_body124_io_Out_67_ready),
    .io_Out_67_valid(bb_for_body124_io_Out_67_valid),
    .io_Out_67_bits_taskID(bb_for_body124_io_Out_67_bits_taskID),
    .io_Out_67_bits_control(bb_for_body124_io_Out_67_bits_control),
    .io_Out_68_ready(bb_for_body124_io_Out_68_ready),
    .io_Out_68_valid(bb_for_body124_io_Out_68_valid),
    .io_Out_68_bits_taskID(bb_for_body124_io_Out_68_bits_taskID),
    .io_Out_68_bits_control(bb_for_body124_io_Out_68_bits_control),
    .io_Out_69_ready(bb_for_body124_io_Out_69_ready),
    .io_Out_69_valid(bb_for_body124_io_Out_69_valid),
    .io_Out_69_bits_taskID(bb_for_body124_io_Out_69_bits_taskID),
    .io_Out_69_bits_control(bb_for_body124_io_Out_69_bits_control),
    .io_Out_70_ready(bb_for_body124_io_Out_70_ready),
    .io_Out_70_valid(bb_for_body124_io_Out_70_valid),
    .io_Out_70_bits_taskID(bb_for_body124_io_Out_70_bits_taskID),
    .io_Out_71_ready(bb_for_body124_io_Out_71_ready),
    .io_Out_71_valid(bb_for_body124_io_Out_71_valid),
    .io_Out_71_bits_taskID(bb_for_body124_io_Out_71_bits_taskID),
    .io_Out_71_bits_control(bb_for_body124_io_Out_71_bits_control),
    .io_Out_72_ready(bb_for_body124_io_Out_72_ready),
    .io_Out_72_valid(bb_for_body124_io_Out_72_valid),
    .io_Out_72_bits_taskID(bb_for_body124_io_Out_72_bits_taskID),
    .io_Out_72_bits_control(bb_for_body124_io_Out_72_bits_control),
    .io_Out_73_ready(bb_for_body124_io_Out_73_ready),
    .io_Out_73_valid(bb_for_body124_io_Out_73_valid),
    .io_Out_73_bits_taskID(bb_for_body124_io_Out_73_bits_taskID),
    .io_Out_73_bits_control(bb_for_body124_io_Out_73_bits_control),
    .io_Out_74_ready(bb_for_body124_io_Out_74_ready),
    .io_Out_74_valid(bb_for_body124_io_Out_74_valid),
    .io_Out_74_bits_taskID(bb_for_body124_io_Out_74_bits_taskID),
    .io_Out_74_bits_control(bb_for_body124_io_Out_74_bits_control),
    .io_Out_75_ready(bb_for_body124_io_Out_75_ready),
    .io_Out_75_valid(bb_for_body124_io_Out_75_valid),
    .io_Out_75_bits_taskID(bb_for_body124_io_Out_75_bits_taskID),
    .io_Out_75_bits_control(bb_for_body124_io_Out_75_bits_control),
    .io_Out_76_ready(bb_for_body124_io_Out_76_ready),
    .io_Out_76_valid(bb_for_body124_io_Out_76_valid),
    .io_Out_76_bits_taskID(bb_for_body124_io_Out_76_bits_taskID),
    .io_Out_76_bits_control(bb_for_body124_io_Out_76_bits_control),
    .io_Out_77_ready(bb_for_body124_io_Out_77_ready),
    .io_Out_77_valid(bb_for_body124_io_Out_77_valid),
    .io_Out_77_bits_taskID(bb_for_body124_io_Out_77_bits_taskID),
    .io_Out_77_bits_control(bb_for_body124_io_Out_77_bits_control),
    .io_Out_78_ready(bb_for_body124_io_Out_78_ready),
    .io_Out_78_valid(bb_for_body124_io_Out_78_valid),
    .io_Out_78_bits_taskID(bb_for_body124_io_Out_78_bits_taskID),
    .io_Out_79_ready(bb_for_body124_io_Out_79_ready),
    .io_Out_79_valid(bb_for_body124_io_Out_79_valid),
    .io_Out_79_bits_taskID(bb_for_body124_io_Out_79_bits_taskID),
    .io_Out_79_bits_control(bb_for_body124_io_Out_79_bits_control),
    .io_Out_80_ready(bb_for_body124_io_Out_80_ready),
    .io_Out_80_valid(bb_for_body124_io_Out_80_valid),
    .io_Out_80_bits_taskID(bb_for_body124_io_Out_80_bits_taskID),
    .io_Out_80_bits_control(bb_for_body124_io_Out_80_bits_control),
    .io_Out_81_ready(bb_for_body124_io_Out_81_ready),
    .io_Out_81_valid(bb_for_body124_io_Out_81_valid),
    .io_Out_81_bits_taskID(bb_for_body124_io_Out_81_bits_taskID),
    .io_Out_81_bits_control(bb_for_body124_io_Out_81_bits_control),
    .io_Out_82_ready(bb_for_body124_io_Out_82_ready),
    .io_Out_82_valid(bb_for_body124_io_Out_82_valid),
    .io_Out_82_bits_taskID(bb_for_body124_io_Out_82_bits_taskID),
    .io_Out_82_bits_control(bb_for_body124_io_Out_82_bits_control),
    .io_Out_83_ready(bb_for_body124_io_Out_83_ready),
    .io_Out_83_valid(bb_for_body124_io_Out_83_valid),
    .io_Out_83_bits_taskID(bb_for_body124_io_Out_83_bits_taskID),
    .io_Out_83_bits_control(bb_for_body124_io_Out_83_bits_control),
    .io_Out_84_ready(bb_for_body124_io_Out_84_ready),
    .io_Out_84_valid(bb_for_body124_io_Out_84_valid),
    .io_Out_84_bits_taskID(bb_for_body124_io_Out_84_bits_taskID),
    .io_Out_84_bits_control(bb_for_body124_io_Out_84_bits_control),
    .io_Out_85_ready(bb_for_body124_io_Out_85_ready),
    .io_Out_85_valid(bb_for_body124_io_Out_85_valid),
    .io_Out_85_bits_taskID(bb_for_body124_io_Out_85_bits_taskID),
    .io_Out_85_bits_control(bb_for_body124_io_Out_85_bits_control),
    .io_Out_86_ready(bb_for_body124_io_Out_86_ready),
    .io_Out_86_valid(bb_for_body124_io_Out_86_valid),
    .io_Out_86_bits_taskID(bb_for_body124_io_Out_86_bits_taskID),
    .io_Out_87_ready(bb_for_body124_io_Out_87_ready),
    .io_Out_87_valid(bb_for_body124_io_Out_87_valid),
    .io_Out_87_bits_taskID(bb_for_body124_io_Out_87_bits_taskID),
    .io_Out_87_bits_control(bb_for_body124_io_Out_87_bits_control),
    .io_Out_88_ready(bb_for_body124_io_Out_88_ready),
    .io_Out_88_valid(bb_for_body124_io_Out_88_valid),
    .io_Out_88_bits_taskID(bb_for_body124_io_Out_88_bits_taskID),
    .io_Out_88_bits_control(bb_for_body124_io_Out_88_bits_control),
    .io_Out_89_ready(bb_for_body124_io_Out_89_ready),
    .io_Out_89_valid(bb_for_body124_io_Out_89_valid),
    .io_Out_89_bits_taskID(bb_for_body124_io_Out_89_bits_taskID),
    .io_Out_89_bits_control(bb_for_body124_io_Out_89_bits_control),
    .io_Out_90_ready(bb_for_body124_io_Out_90_ready),
    .io_Out_90_valid(bb_for_body124_io_Out_90_valid),
    .io_Out_90_bits_taskID(bb_for_body124_io_Out_90_bits_taskID),
    .io_Out_90_bits_control(bb_for_body124_io_Out_90_bits_control),
    .io_Out_91_ready(bb_for_body124_io_Out_91_ready),
    .io_Out_91_valid(bb_for_body124_io_Out_91_valid),
    .io_Out_91_bits_taskID(bb_for_body124_io_Out_91_bits_taskID),
    .io_Out_91_bits_control(bb_for_body124_io_Out_91_bits_control),
    .io_Out_92_ready(bb_for_body124_io_Out_92_ready),
    .io_Out_92_valid(bb_for_body124_io_Out_92_valid),
    .io_Out_92_bits_taskID(bb_for_body124_io_Out_92_bits_taskID),
    .io_Out_92_bits_control(bb_for_body124_io_Out_92_bits_control),
    .io_predicateIn_0_ready(bb_for_body124_io_predicateIn_0_ready),
    .io_predicateIn_0_valid(bb_for_body124_io_predicateIn_0_valid),
    .io_predicateIn_0_bits_taskID(bb_for_body124_io_predicateIn_0_bits_taskID),
    .io_predicateIn_0_bits_control(bb_for_body124_io_predicateIn_0_bits_control),
    .io_predicateIn_1_ready(bb_for_body124_io_predicateIn_1_ready),
    .io_predicateIn_1_valid(bb_for_body124_io_predicateIn_1_valid),
    .io_predicateIn_1_bits_taskID(bb_for_body124_io_predicateIn_1_bits_taskID),
    .io_predicateIn_1_bits_control(bb_for_body124_io_predicateIn_1_bits_control)
  );
  ComputeNode binaryOp_mul0 ( // @[extracted_function_conv.scala 89:29]
    .clock(binaryOp_mul0_clock),
    .reset(binaryOp_mul0_reset),
    .io_enable_ready(binaryOp_mul0_io_enable_ready),
    .io_enable_valid(binaryOp_mul0_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul0_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul0_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul0_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul0_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul0_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul0_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul0_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul0_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul0_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul0_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul0_io_RightIO_bits_data)
  );
  ComputeNode_1 binaryOp_add1 ( // @[extracted_function_conv.scala 92:29]
    .clock(binaryOp_add1_clock),
    .reset(binaryOp_add1_reset),
    .io_enable_ready(binaryOp_add1_io_enable_ready),
    .io_enable_valid(binaryOp_add1_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add1_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add1_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add1_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add1_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add1_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add1_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add1_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add1_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add1_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add1_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add1_io_RightIO_bits_data)
  );
  GepNode Gep_arrayidx252 ( // @[extracted_function_conv.scala 95:31]
    .clock(Gep_arrayidx252_clock),
    .reset(Gep_arrayidx252_reset),
    .io_enable_ready(Gep_arrayidx252_io_enable_ready),
    .io_enable_valid(Gep_arrayidx252_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx252_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx252_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx252_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx252_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx252_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx252_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx252_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx252_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx252_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx252_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx252_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx252_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx252_io_idx_0_valid)
  );
  GepNode_1 Gep_arrayidx383 ( // @[extracted_function_conv.scala 98:31]
    .clock(Gep_arrayidx383_clock),
    .reset(Gep_arrayidx383_reset),
    .io_enable_ready(Gep_arrayidx383_io_enable_ready),
    .io_enable_valid(Gep_arrayidx383_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx383_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx383_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx383_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx383_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx383_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx383_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx383_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx383_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx383_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx383_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx383_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx383_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx383_io_idx_0_valid)
  );
  GepNode_2 Gep_arrayidx514 ( // @[extracted_function_conv.scala 101:31]
    .clock(Gep_arrayidx514_clock),
    .reset(Gep_arrayidx514_reset),
    .io_enable_ready(Gep_arrayidx514_io_enable_ready),
    .io_enable_valid(Gep_arrayidx514_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx514_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx514_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx514_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx514_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx514_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx514_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx514_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx514_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx514_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx514_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx514_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx514_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx514_io_idx_0_valid)
  );
  GepNode_3 Gep_arrayidx625 ( // @[extracted_function_conv.scala 104:31]
    .clock(Gep_arrayidx625_clock),
    .reset(Gep_arrayidx625_reset),
    .io_enable_ready(Gep_arrayidx625_io_enable_ready),
    .io_enable_valid(Gep_arrayidx625_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx625_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx625_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx625_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx625_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx625_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx625_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx625_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx625_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx625_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx625_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx625_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx625_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx625_io_idx_0_valid)
  );
  GepNode_4 Gep_arrayidx746 ( // @[extracted_function_conv.scala 107:31]
    .clock(Gep_arrayidx746_clock),
    .reset(Gep_arrayidx746_reset),
    .io_enable_ready(Gep_arrayidx746_io_enable_ready),
    .io_enable_valid(Gep_arrayidx746_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx746_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx746_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx746_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx746_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx746_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx746_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx746_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx746_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx746_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx746_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx746_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx746_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx746_io_idx_0_valid)
  );
  GepNode_5 Gep_arrayidx867 ( // @[extracted_function_conv.scala 110:31]
    .clock(Gep_arrayidx867_clock),
    .reset(Gep_arrayidx867_reset),
    .io_enable_ready(Gep_arrayidx867_io_enable_ready),
    .io_enable_valid(Gep_arrayidx867_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx867_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx867_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx867_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx867_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx867_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx867_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx867_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx867_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx867_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx867_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx867_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx867_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx867_io_idx_0_valid)
  );
  GepNode_6 Gep_arrayidx978 ( // @[extracted_function_conv.scala 113:31]
    .clock(Gep_arrayidx978_clock),
    .reset(Gep_arrayidx978_reset),
    .io_enable_ready(Gep_arrayidx978_io_enable_ready),
    .io_enable_valid(Gep_arrayidx978_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx978_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx978_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx978_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx978_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx978_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx978_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx978_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx978_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx978_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx978_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx978_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx978_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx978_io_idx_0_valid)
  );
  GepNode_7 Gep_arrayidx1099 ( // @[extracted_function_conv.scala 116:32]
    .clock(Gep_arrayidx1099_clock),
    .reset(Gep_arrayidx1099_reset),
    .io_enable_ready(Gep_arrayidx1099_io_enable_ready),
    .io_enable_valid(Gep_arrayidx1099_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx1099_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx1099_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx1099_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx1099_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx1099_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx1099_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx1099_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx1099_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx1099_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx1099_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx1099_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx1099_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx1099_io_idx_0_valid)
  );
  UBranchNode br_10 ( // @[extracted_function_conv.scala 119:21]
    .clock(br_10_clock),
    .reset(br_10_reset),
    .io_enable_ready(br_10_io_enable_ready),
    .io_enable_valid(br_10_io_enable_valid),
    .io_enable_bits_taskID(br_10_io_enable_bits_taskID),
    .io_enable_bits_control(br_10_io_enable_bits_control),
    .io_Out_0_ready(br_10_io_Out_0_ready),
    .io_Out_0_valid(br_10_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_10_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_10_io_Out_0_bits_control)
  );
  RetNode2 ret_11 ( // @[extracted_function_conv.scala 122:22]
    .clock(ret_11_clock),
    .reset(ret_11_reset),
    .io_In_enable_ready(ret_11_io_In_enable_ready),
    .io_In_enable_valid(ret_11_io_In_enable_valid),
    .io_In_enable_bits_taskID(ret_11_io_In_enable_bits_taskID),
    .io_In_enable_bits_control(ret_11_io_In_enable_bits_control),
    .io_Out_ready(ret_11_io_Out_ready),
    .io_Out_valid(ret_11_io_Out_valid),
    .io_Out_bits_enable_taskID(ret_11_io_Out_bits_enable_taskID),
    .io_Out_bits_enable_control(ret_11_io_Out_bits_enable_control)
  );
  PhiFastNode phi_conv_s1_y_031312 ( // @[extracted_function_conv.scala 125:36]
    .clock(phi_conv_s1_y_031312_clock),
    .reset(phi_conv_s1_y_031312_reset),
    .io_enable_ready(phi_conv_s1_y_031312_io_enable_ready),
    .io_enable_valid(phi_conv_s1_y_031312_io_enable_valid),
    .io_enable_bits_control(phi_conv_s1_y_031312_io_enable_bits_control),
    .io_InData_0_ready(phi_conv_s1_y_031312_io_InData_0_ready),
    .io_InData_0_valid(phi_conv_s1_y_031312_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_conv_s1_y_031312_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi_conv_s1_y_031312_io_InData_1_ready),
    .io_InData_1_valid(phi_conv_s1_y_031312_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_conv_s1_y_031312_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_conv_s1_y_031312_io_InData_1_bits_data),
    .io_Mask_ready(phi_conv_s1_y_031312_io_Mask_ready),
    .io_Mask_valid(phi_conv_s1_y_031312_io_Mask_valid),
    .io_Mask_bits(phi_conv_s1_y_031312_io_Mask_bits),
    .io_Out_0_ready(phi_conv_s1_y_031312_io_Out_0_ready),
    .io_Out_0_valid(phi_conv_s1_y_031312_io_Out_0_valid),
    .io_Out_0_bits_data(phi_conv_s1_y_031312_io_Out_0_bits_data),
    .io_Out_1_ready(phi_conv_s1_y_031312_io_Out_1_ready),
    .io_Out_1_valid(phi_conv_s1_y_031312_io_Out_1_valid),
    .io_Out_1_bits_data(phi_conv_s1_y_031312_io_Out_1_bits_data),
    .io_Out_2_ready(phi_conv_s1_y_031312_io_Out_2_ready),
    .io_Out_2_valid(phi_conv_s1_y_031312_io_Out_2_valid),
    .io_Out_2_bits_data(phi_conv_s1_y_031312_io_Out_2_bits_data),
    .io_Out_3_ready(phi_conv_s1_y_031312_io_Out_3_ready),
    .io_Out_3_valid(phi_conv_s1_y_031312_io_Out_3_valid),
    .io_Out_3_bits_data(phi_conv_s1_y_031312_io_Out_3_bits_data)
  );
  ComputeNode_2 binaryOp_mul113 ( // @[extracted_function_conv.scala 128:31]
    .clock(binaryOp_mul113_clock),
    .reset(binaryOp_mul113_reset),
    .io_enable_ready(binaryOp_mul113_io_enable_ready),
    .io_enable_valid(binaryOp_mul113_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul113_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul113_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul113_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul113_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul113_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_mul113_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_mul113_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_mul113_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_mul113_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul113_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul113_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul113_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul113_io_RightIO_valid)
  );
  ComputeNode_3 binaryOp_add214 ( // @[extracted_function_conv.scala 131:31]
    .clock(binaryOp_add214_clock),
    .reset(binaryOp_add214_reset),
    .io_enable_ready(binaryOp_add214_io_enable_ready),
    .io_enable_valid(binaryOp_add214_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add214_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add214_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add214_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add214_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add214_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add214_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add214_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add214_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add214_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add214_io_RightIO_valid)
  );
  ComputeNode_4 binaryOp_mul315 ( // @[extracted_function_conv.scala 134:31]
    .clock(binaryOp_mul315_clock),
    .reset(binaryOp_mul315_reset),
    .io_enable_ready(binaryOp_mul315_io_enable_ready),
    .io_enable_valid(binaryOp_mul315_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul315_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul315_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul315_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul315_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul315_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul315_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul315_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul315_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul315_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul315_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul315_io_RightIO_bits_data)
  );
  ComputeNode_5 binaryOp_sub16 ( // @[extracted_function_conv.scala 137:30]
    .clock(binaryOp_sub16_clock),
    .reset(binaryOp_sub16_reset),
    .io_enable_ready(binaryOp_sub16_io_enable_ready),
    .io_enable_valid(binaryOp_sub16_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_sub16_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_sub16_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_sub16_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_sub16_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_sub16_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_sub16_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_sub16_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_sub16_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_sub16_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_sub16_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_sub16_io_RightIO_bits_data)
  );
  ComputeNode_6 binaryOp_add417 ( // @[extracted_function_conv.scala 140:31]
    .clock(binaryOp_add417_clock),
    .reset(binaryOp_add417_reset),
    .io_enable_ready(binaryOp_add417_io_enable_ready),
    .io_enable_valid(binaryOp_add417_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add417_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add417_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add417_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add417_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add417_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add417_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add417_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add417_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add417_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add417_io_RightIO_valid)
  );
  ComputeNode_7 binaryOp_mul518 ( // @[extracted_function_conv.scala 143:31]
    .clock(binaryOp_mul518_clock),
    .reset(binaryOp_mul518_reset),
    .io_enable_ready(binaryOp_mul518_io_enable_ready),
    .io_enable_valid(binaryOp_mul518_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul518_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul518_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul518_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul518_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul518_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul518_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul518_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul518_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul518_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul518_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul518_io_RightIO_bits_data)
  );
  ComputeNode_8 binaryOp_sub619 ( // @[extracted_function_conv.scala 146:31]
    .clock(binaryOp_sub619_clock),
    .reset(binaryOp_sub619_reset),
    .io_enable_ready(binaryOp_sub619_io_enable_ready),
    .io_enable_valid(binaryOp_sub619_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_sub619_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_sub619_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_sub619_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_sub619_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_sub619_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_sub619_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_sub619_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_sub619_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_sub619_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_sub619_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_sub619_io_RightIO_bits_data)
  );
  ComputeNode_9 binaryOp_mul720 ( // @[extracted_function_conv.scala 149:31]
    .clock(binaryOp_mul720_clock),
    .reset(binaryOp_mul720_reset),
    .io_enable_ready(binaryOp_mul720_io_enable_ready),
    .io_enable_valid(binaryOp_mul720_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul720_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul720_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul720_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul720_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul720_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul720_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul720_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul720_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul720_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul720_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul720_io_RightIO_bits_data)
  );
  ComputeNode_10 binaryOp_mul821 ( // @[extracted_function_conv.scala 152:31]
    .clock(binaryOp_mul821_clock),
    .reset(binaryOp_mul821_reset),
    .io_enable_ready(binaryOp_mul821_io_enable_ready),
    .io_enable_valid(binaryOp_mul821_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul821_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul821_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul821_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul821_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul821_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul821_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul821_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul821_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul821_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul821_io_RightIO_valid)
  );
  UBranchNode_1 br_22 ( // @[extracted_function_conv.scala 155:21]
    .clock(br_22_clock),
    .reset(br_22_reset),
    .io_enable_ready(br_22_io_enable_ready),
    .io_enable_valid(br_22_io_enable_valid),
    .io_enable_bits_taskID(br_22_io_enable_bits_taskID),
    .io_enable_bits_control(br_22_io_enable_bits_control),
    .io_Out_0_ready(br_22_io_Out_0_ready),
    .io_Out_0_valid(br_22_io_Out_0_valid),
    .io_Out_0_bits_taskID(br_22_io_Out_0_bits_taskID),
    .io_Out_0_bits_control(br_22_io_Out_0_bits_control)
  );
  ComputeNode_11 binaryOp_inc12023 ( // @[extracted_function_conv.scala 158:33]
    .clock(binaryOp_inc12023_clock),
    .reset(binaryOp_inc12023_reset),
    .io_enable_ready(binaryOp_inc12023_io_enable_ready),
    .io_enable_valid(binaryOp_inc12023_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_inc12023_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_inc12023_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_inc12023_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_inc12023_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_inc12023_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_inc12023_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_inc12023_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_inc12023_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_inc12023_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_inc12023_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_inc12023_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_inc12023_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_inc12023_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_inc12023_io_RightIO_valid)
  );
  ComputeNode_12 icmp_exitcond31424 ( // @[extracted_function_conv.scala 161:34]
    .clock(icmp_exitcond31424_clock),
    .reset(icmp_exitcond31424_reset),
    .io_enable_ready(icmp_exitcond31424_io_enable_ready),
    .io_enable_valid(icmp_exitcond31424_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond31424_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond31424_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond31424_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond31424_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond31424_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond31424_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond31424_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond31424_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond31424_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond31424_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond31424_io_RightIO_valid)
  );
  CBranchNodeVariable br_25 ( // @[extracted_function_conv.scala 164:21]
    .clock(br_25_clock),
    .reset(br_25_reset),
    .io_enable_ready(br_25_io_enable_ready),
    .io_enable_valid(br_25_io_enable_valid),
    .io_enable_bits_taskID(br_25_io_enable_bits_taskID),
    .io_enable_bits_control(br_25_io_enable_bits_control),
    .io_CmpIO_ready(br_25_io_CmpIO_ready),
    .io_CmpIO_valid(br_25_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_25_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_25_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_25_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_25_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_25_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_25_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_25_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_25_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_25_io_FalseOutput_0_bits_control)
  );
  PhiFastNode_1 phi_conv_s1_x_031226 ( // @[extracted_function_conv.scala 167:36]
    .clock(phi_conv_s1_x_031226_clock),
    .reset(phi_conv_s1_x_031226_reset),
    .io_enable_ready(phi_conv_s1_x_031226_io_enable_ready),
    .io_enable_valid(phi_conv_s1_x_031226_io_enable_valid),
    .io_enable_bits_control(phi_conv_s1_x_031226_io_enable_bits_control),
    .io_InData_0_ready(phi_conv_s1_x_031226_io_InData_0_ready),
    .io_InData_0_valid(phi_conv_s1_x_031226_io_InData_0_valid),
    .io_InData_0_bits_taskID(phi_conv_s1_x_031226_io_InData_0_bits_taskID),
    .io_InData_1_ready(phi_conv_s1_x_031226_io_InData_1_ready),
    .io_InData_1_valid(phi_conv_s1_x_031226_io_InData_1_valid),
    .io_InData_1_bits_taskID(phi_conv_s1_x_031226_io_InData_1_bits_taskID),
    .io_InData_1_bits_data(phi_conv_s1_x_031226_io_InData_1_bits_data),
    .io_Mask_ready(phi_conv_s1_x_031226_io_Mask_ready),
    .io_Mask_valid(phi_conv_s1_x_031226_io_Mask_valid),
    .io_Mask_bits(phi_conv_s1_x_031226_io_Mask_bits),
    .io_Out_0_ready(phi_conv_s1_x_031226_io_Out_0_ready),
    .io_Out_0_valid(phi_conv_s1_x_031226_io_Out_0_valid),
    .io_Out_0_bits_data(phi_conv_s1_x_031226_io_Out_0_bits_data),
    .io_Out_1_ready(phi_conv_s1_x_031226_io_Out_1_ready),
    .io_Out_1_valid(phi_conv_s1_x_031226_io_Out_1_valid),
    .io_Out_1_bits_data(phi_conv_s1_x_031226_io_Out_1_bits_data),
    .io_Out_2_ready(phi_conv_s1_x_031226_io_Out_2_ready),
    .io_Out_2_valid(phi_conv_s1_x_031226_io_Out_2_valid),
    .io_Out_2_bits_data(phi_conv_s1_x_031226_io_Out_2_bits_data),
    .io_Out_3_ready(phi_conv_s1_x_031226_io_Out_3_ready),
    .io_Out_3_valid(phi_conv_s1_x_031226_io_Out_3_valid),
    .io_Out_3_bits_data(phi_conv_s1_x_031226_io_Out_3_bits_data)
  );
  ComputeNode_13 binaryOp_add1327 ( // @[extracted_function_conv.scala 170:32]
    .clock(binaryOp_add1327_clock),
    .reset(binaryOp_add1327_reset),
    .io_enable_ready(binaryOp_add1327_io_enable_ready),
    .io_enable_valid(binaryOp_add1327_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add1327_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add1327_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add1327_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add1327_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add1327_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add1327_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add1327_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add1327_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add1327_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add1327_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add1327_io_RightIO_bits_data)
  );
  GepNode_8 Gep_arrayidx28 ( // @[extracted_function_conv.scala 173:30]
    .clock(Gep_arrayidx28_clock),
    .reset(Gep_arrayidx28_reset),
    .io_enable_ready(Gep_arrayidx28_io_enable_ready),
    .io_enable_valid(Gep_arrayidx28_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx28_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx28_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx28_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx28_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx28_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx28_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx28_io_Out_0_bits_data),
    .io_Out_1_ready(Gep_arrayidx28_io_Out_1_ready),
    .io_Out_1_valid(Gep_arrayidx28_io_Out_1_valid),
    .io_Out_1_bits_taskID(Gep_arrayidx28_io_Out_1_bits_taskID),
    .io_Out_1_bits_data(Gep_arrayidx28_io_Out_1_bits_data),
    .io_Out_2_ready(Gep_arrayidx28_io_Out_2_ready),
    .io_Out_2_valid(Gep_arrayidx28_io_Out_2_valid),
    .io_Out_2_bits_taskID(Gep_arrayidx28_io_Out_2_bits_taskID),
    .io_Out_2_bits_data(Gep_arrayidx28_io_Out_2_bits_data),
    .io_Out_3_ready(Gep_arrayidx28_io_Out_3_ready),
    .io_Out_3_valid(Gep_arrayidx28_io_Out_3_valid),
    .io_Out_3_bits_taskID(Gep_arrayidx28_io_Out_3_bits_taskID),
    .io_Out_3_bits_data(Gep_arrayidx28_io_Out_3_bits_data),
    .io_Out_4_ready(Gep_arrayidx28_io_Out_4_ready),
    .io_Out_4_valid(Gep_arrayidx28_io_Out_4_valid),
    .io_Out_4_bits_taskID(Gep_arrayidx28_io_Out_4_bits_taskID),
    .io_Out_4_bits_data(Gep_arrayidx28_io_Out_4_bits_data),
    .io_Out_5_ready(Gep_arrayidx28_io_Out_5_ready),
    .io_Out_5_valid(Gep_arrayidx28_io_Out_5_valid),
    .io_Out_5_bits_taskID(Gep_arrayidx28_io_Out_5_bits_taskID),
    .io_Out_5_bits_data(Gep_arrayidx28_io_Out_5_bits_data),
    .io_Out_6_ready(Gep_arrayidx28_io_Out_6_ready),
    .io_Out_6_valid(Gep_arrayidx28_io_Out_6_valid),
    .io_Out_6_bits_taskID(Gep_arrayidx28_io_Out_6_bits_taskID),
    .io_Out_6_bits_data(Gep_arrayidx28_io_Out_6_bits_data),
    .io_Out_7_ready(Gep_arrayidx28_io_Out_7_ready),
    .io_Out_7_valid(Gep_arrayidx28_io_Out_7_valid),
    .io_Out_7_bits_taskID(Gep_arrayidx28_io_Out_7_bits_taskID),
    .io_Out_7_bits_data(Gep_arrayidx28_io_Out_7_bits_data),
    .io_Out_8_ready(Gep_arrayidx28_io_Out_8_ready),
    .io_Out_8_valid(Gep_arrayidx28_io_Out_8_valid),
    .io_Out_8_bits_taskID(Gep_arrayidx28_io_Out_8_bits_taskID),
    .io_Out_8_bits_data(Gep_arrayidx28_io_Out_8_bits_data),
    .io_Out_9_ready(Gep_arrayidx28_io_Out_9_ready),
    .io_Out_9_valid(Gep_arrayidx28_io_Out_9_valid),
    .io_Out_9_bits_taskID(Gep_arrayidx28_io_Out_9_bits_taskID),
    .io_Out_9_bits_data(Gep_arrayidx28_io_Out_9_bits_data),
    .io_baseAddress_ready(Gep_arrayidx28_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx28_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx28_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx28_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx28_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx28_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx28_io_idx_0_bits_data)
  );
  UnTypLoad ld_29 ( // @[extracted_function_conv.scala 176:21]
    .clock(ld_29_clock),
    .reset(ld_29_reset),
    .io_enable_ready(ld_29_io_enable_ready),
    .io_enable_valid(ld_29_io_enable_valid),
    .io_enable_bits_taskID(ld_29_io_enable_bits_taskID),
    .io_enable_bits_control(ld_29_io_enable_bits_control),
    .io_Out_0_ready(ld_29_io_Out_0_ready),
    .io_Out_0_valid(ld_29_io_Out_0_valid),
    .io_Out_0_bits_data(ld_29_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_29_io_GepAddr_ready),
    .io_GepAddr_valid(ld_29_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_29_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_29_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_29_io_GepAddr_bits_data),
    .io_memReq_ready(ld_29_io_memReq_ready),
    .io_memReq_valid(ld_29_io_memReq_valid),
    .io_memReq_bits_address(ld_29_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_29_io_memReq_bits_taskID),
    .io_memResp_valid(ld_29_io_memResp_valid),
    .io_memResp_data(ld_29_io_memResp_data)
  );
  UnTypLoad_1 ld_30 ( // @[extracted_function_conv.scala 179:21]
    .clock(ld_30_clock),
    .reset(ld_30_reset),
    .io_enable_ready(ld_30_io_enable_ready),
    .io_enable_valid(ld_30_io_enable_valid),
    .io_enable_bits_taskID(ld_30_io_enable_bits_taskID),
    .io_enable_bits_control(ld_30_io_enable_bits_control),
    .io_Out_0_ready(ld_30_io_Out_0_ready),
    .io_Out_0_valid(ld_30_io_Out_0_valid),
    .io_Out_0_bits_data(ld_30_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_30_io_GepAddr_ready),
    .io_GepAddr_valid(ld_30_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_30_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_30_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_30_io_GepAddr_bits_data),
    .io_memReq_ready(ld_30_io_memReq_ready),
    .io_memReq_valid(ld_30_io_memReq_valid),
    .io_memReq_bits_address(ld_30_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_30_io_memReq_bits_taskID),
    .io_memResp_valid(ld_30_io_memResp_valid),
    .io_memResp_data(ld_30_io_memResp_data)
  );
  ComputeNode_14 binaryOp_add1531 ( // @[extracted_function_conv.scala 182:32]
    .clock(binaryOp_add1531_clock),
    .reset(binaryOp_add1531_reset),
    .io_enable_ready(binaryOp_add1531_io_enable_ready),
    .io_enable_valid(binaryOp_add1531_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add1531_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add1531_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add1531_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add1531_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add1531_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add1531_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add1531_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add1531_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add1531_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add1531_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add1531_io_RightIO_bits_data)
  );
  ComputeNode_15 binaryOp_mul1632 ( // @[extracted_function_conv.scala 185:32]
    .clock(binaryOp_mul1632_clock),
    .reset(binaryOp_mul1632_reset),
    .io_enable_ready(binaryOp_mul1632_io_enable_ready),
    .io_enable_valid(binaryOp_mul1632_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul1632_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul1632_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul1632_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul1632_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul1632_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul1632_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul1632_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul1632_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul1632_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul1632_io_RightIO_valid)
  );
  ComputeNode_16 binaryOp_sub1733 ( // @[extracted_function_conv.scala 188:32]
    .clock(binaryOp_sub1733_clock),
    .reset(binaryOp_sub1733_reset),
    .io_enable_ready(binaryOp_sub1733_io_enable_ready),
    .io_enable_valid(binaryOp_sub1733_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_sub1733_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_sub1733_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_sub1733_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_sub1733_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_sub1733_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_sub1733_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_sub1733_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_sub1733_io_Out_1_bits_data),
    .io_Out_2_ready(binaryOp_sub1733_io_Out_2_ready),
    .io_Out_2_valid(binaryOp_sub1733_io_Out_2_valid),
    .io_Out_2_bits_data(binaryOp_sub1733_io_Out_2_bits_data),
    .io_LeftIO_ready(binaryOp_sub1733_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_sub1733_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_sub1733_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_sub1733_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_sub1733_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_sub1733_io_RightIO_bits_data)
  );
  GepNode_9 Gep_arrayidx1834 ( // @[extracted_function_conv.scala 191:32]
    .clock(Gep_arrayidx1834_clock),
    .reset(Gep_arrayidx1834_reset),
    .io_enable_ready(Gep_arrayidx1834_io_enable_ready),
    .io_enable_valid(Gep_arrayidx1834_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx1834_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx1834_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx1834_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx1834_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx1834_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx1834_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx1834_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx1834_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx1834_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx1834_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx1834_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx1834_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx1834_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx1834_io_idx_0_bits_data)
  );
  UnTypLoad_2 ld_35 ( // @[extracted_function_conv.scala 194:21]
    .clock(ld_35_clock),
    .reset(ld_35_reset),
    .io_enable_ready(ld_35_io_enable_ready),
    .io_enable_valid(ld_35_io_enable_valid),
    .io_enable_bits_taskID(ld_35_io_enable_bits_taskID),
    .io_enable_bits_control(ld_35_io_enable_bits_control),
    .io_Out_0_ready(ld_35_io_Out_0_ready),
    .io_Out_0_valid(ld_35_io_Out_0_valid),
    .io_Out_0_bits_data(ld_35_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_35_io_GepAddr_ready),
    .io_GepAddr_valid(ld_35_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_35_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_35_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_35_io_GepAddr_bits_data),
    .io_memReq_ready(ld_35_io_memReq_ready),
    .io_memReq_valid(ld_35_io_memReq_valid),
    .io_memReq_bits_address(ld_35_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_35_io_memReq_bits_taskID),
    .io_memResp_valid(ld_35_io_memResp_valid),
    .io_memResp_data(ld_35_io_memResp_data)
  );
  ZextNode sextconv1936 ( // @[extracted_function_conv.scala 197:28]
    .clock(sextconv1936_clock),
    .reset(sextconv1936_reset),
    .io_Input_ready(sextconv1936_io_Input_ready),
    .io_Input_valid(sextconv1936_io_Input_valid),
    .io_Input_bits_data(sextconv1936_io_Input_bits_data),
    .io_enable_ready(sextconv1936_io_enable_ready),
    .io_enable_valid(sextconv1936_io_enable_valid),
    .io_enable_bits_taskID(sextconv1936_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv1936_io_Out_0_ready),
    .io_Out_0_valid(sextconv1936_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv1936_io_Out_0_bits_data)
  );
  ComputeNode_17 binaryOp_mul2037 ( // @[extracted_function_conv.scala 200:32]
    .clock(binaryOp_mul2037_clock),
    .reset(binaryOp_mul2037_reset),
    .io_enable_ready(binaryOp_mul2037_io_enable_ready),
    .io_enable_valid(binaryOp_mul2037_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul2037_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul2037_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul2037_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul2037_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul2037_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul2037_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul2037_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul2037_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul2037_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul2037_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul2037_io_RightIO_bits_data)
  );
  ComputeNode_18 binaryOp_add2138 ( // @[extracted_function_conv.scala 203:32]
    .clock(binaryOp_add2138_clock),
    .reset(binaryOp_add2138_reset),
    .io_enable_ready(binaryOp_add2138_io_enable_ready),
    .io_enable_valid(binaryOp_add2138_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add2138_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add2138_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add2138_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add2138_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add2138_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add2138_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add2138_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add2138_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add2138_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add2138_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add2138_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add2138_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add2138_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add2138_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add2138_io_RightIO_bits_data)
  );
  UnTypStore st_39 ( // @[extracted_function_conv.scala 206:21]
    .clock(st_39_clock),
    .reset(st_39_reset),
    .io_enable_ready(st_39_io_enable_ready),
    .io_enable_valid(st_39_io_enable_valid),
    .io_enable_bits_taskID(st_39_io_enable_bits_taskID),
    .io_enable_bits_control(st_39_io_enable_bits_control),
    .io_GepAddr_ready(st_39_io_GepAddr_ready),
    .io_GepAddr_valid(st_39_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_39_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_39_io_GepAddr_bits_data),
    .io_inData_ready(st_39_io_inData_ready),
    .io_inData_valid(st_39_io_inData_valid),
    .io_inData_bits_taskID(st_39_io_inData_bits_taskID),
    .io_inData_bits_data(st_39_io_inData_bits_data),
    .io_memReq_ready(st_39_io_memReq_ready),
    .io_memReq_valid(st_39_io_memReq_valid),
    .io_memReq_bits_address(st_39_io_memReq_bits_address),
    .io_memReq_bits_data(st_39_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_39_io_memReq_bits_taskID),
    .io_memResp_valid(st_39_io_memResp_valid)
  );
  UnTypLoad_3 ld_40 ( // @[extracted_function_conv.scala 209:21]
    .clock(ld_40_clock),
    .reset(ld_40_reset),
    .io_enable_ready(ld_40_io_enable_ready),
    .io_enable_valid(ld_40_io_enable_valid),
    .io_enable_bits_taskID(ld_40_io_enable_bits_taskID),
    .io_enable_bits_control(ld_40_io_enable_bits_control),
    .io_Out_0_ready(ld_40_io_Out_0_ready),
    .io_Out_0_valid(ld_40_io_Out_0_valid),
    .io_Out_0_bits_data(ld_40_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_40_io_GepAddr_ready),
    .io_GepAddr_valid(ld_40_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_40_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_40_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_40_io_GepAddr_bits_data),
    .io_memReq_ready(ld_40_io_memReq_ready),
    .io_memReq_valid(ld_40_io_memReq_valid),
    .io_memReq_bits_address(ld_40_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_40_io_memReq_bits_taskID),
    .io_memResp_valid(ld_40_io_memResp_valid),
    .io_memResp_data(ld_40_io_memResp_data)
  );
  ComputeNode_19 binaryOp_add2941 ( // @[extracted_function_conv.scala 212:32]
    .clock(binaryOp_add2941_clock),
    .reset(binaryOp_add2941_reset),
    .io_enable_ready(binaryOp_add2941_io_enable_ready),
    .io_enable_valid(binaryOp_add2941_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add2941_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add2941_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add2941_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add2941_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add2941_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add2941_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add2941_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add2941_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add2941_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add2941_io_RightIO_valid)
  );
  GepNode_10 Gep_arrayidx3042 ( // @[extracted_function_conv.scala 215:32]
    .clock(Gep_arrayidx3042_clock),
    .reset(Gep_arrayidx3042_reset),
    .io_enable_ready(Gep_arrayidx3042_io_enable_ready),
    .io_enable_valid(Gep_arrayidx3042_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx3042_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx3042_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx3042_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx3042_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx3042_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx3042_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx3042_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx3042_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx3042_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx3042_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx3042_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx3042_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx3042_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx3042_io_idx_0_bits_data)
  );
  UnTypLoad_4 ld_43 ( // @[extracted_function_conv.scala 218:21]
    .clock(ld_43_clock),
    .reset(ld_43_reset),
    .io_enable_ready(ld_43_io_enable_ready),
    .io_enable_valid(ld_43_io_enable_valid),
    .io_enable_bits_taskID(ld_43_io_enable_bits_taskID),
    .io_enable_bits_control(ld_43_io_enable_bits_control),
    .io_Out_0_ready(ld_43_io_Out_0_ready),
    .io_Out_0_valid(ld_43_io_Out_0_valid),
    .io_Out_0_bits_data(ld_43_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_43_io_GepAddr_ready),
    .io_GepAddr_valid(ld_43_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_43_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_43_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_43_io_GepAddr_bits_data),
    .io_memReq_ready(ld_43_io_memReq_ready),
    .io_memReq_valid(ld_43_io_memReq_valid),
    .io_memReq_bits_address(ld_43_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_43_io_memReq_bits_taskID),
    .io_memResp_valid(ld_43_io_memResp_valid),
    .io_memResp_data(ld_43_io_memResp_data)
  );
  ZextNode_1 sextconv3244 ( // @[extracted_function_conv.scala 221:28]
    .clock(sextconv3244_clock),
    .reset(sextconv3244_reset),
    .io_Input_ready(sextconv3244_io_Input_ready),
    .io_Input_valid(sextconv3244_io_Input_valid),
    .io_Input_bits_data(sextconv3244_io_Input_bits_data),
    .io_enable_ready(sextconv3244_io_enable_ready),
    .io_enable_valid(sextconv3244_io_enable_valid),
    .io_enable_bits_taskID(sextconv3244_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv3244_io_Out_0_ready),
    .io_Out_0_valid(sextconv3244_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv3244_io_Out_0_bits_data)
  );
  ComputeNode_20 binaryOp_mul3345 ( // @[extracted_function_conv.scala 224:32]
    .clock(binaryOp_mul3345_clock),
    .reset(binaryOp_mul3345_reset),
    .io_enable_ready(binaryOp_mul3345_io_enable_ready),
    .io_enable_valid(binaryOp_mul3345_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul3345_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul3345_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul3345_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul3345_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul3345_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul3345_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul3345_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul3345_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul3345_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul3345_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul3345_io_RightIO_bits_data)
  );
  ComputeNode_21 binaryOp_add3446 ( // @[extracted_function_conv.scala 227:32]
    .clock(binaryOp_add3446_clock),
    .reset(binaryOp_add3446_reset),
    .io_enable_ready(binaryOp_add3446_io_enable_ready),
    .io_enable_valid(binaryOp_add3446_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add3446_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add3446_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add3446_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add3446_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add3446_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add3446_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add3446_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add3446_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add3446_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add3446_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add3446_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add3446_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add3446_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add3446_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add3446_io_RightIO_bits_data)
  );
  UnTypStore_1 st_47 ( // @[extracted_function_conv.scala 230:21]
    .clock(st_47_clock),
    .reset(st_47_reset),
    .io_enable_ready(st_47_io_enable_ready),
    .io_enable_valid(st_47_io_enable_valid),
    .io_enable_bits_taskID(st_47_io_enable_bits_taskID),
    .io_enable_bits_control(st_47_io_enable_bits_control),
    .io_GepAddr_ready(st_47_io_GepAddr_ready),
    .io_GepAddr_valid(st_47_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_47_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_47_io_GepAddr_bits_data),
    .io_inData_ready(st_47_io_inData_ready),
    .io_inData_valid(st_47_io_inData_valid),
    .io_inData_bits_taskID(st_47_io_inData_bits_taskID),
    .io_inData_bits_data(st_47_io_inData_bits_data),
    .io_memReq_ready(st_47_io_memReq_ready),
    .io_memReq_valid(st_47_io_memReq_valid),
    .io_memReq_bits_address(st_47_io_memReq_bits_address),
    .io_memReq_bits_data(st_47_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_47_io_memReq_bits_taskID),
    .io_memResp_valid(st_47_io_memResp_valid)
  );
  UnTypLoad_5 ld_48 ( // @[extracted_function_conv.scala 233:21]
    .clock(ld_48_clock),
    .reset(ld_48_reset),
    .io_enable_ready(ld_48_io_enable_ready),
    .io_enable_valid(ld_48_io_enable_valid),
    .io_enable_bits_taskID(ld_48_io_enable_bits_taskID),
    .io_enable_bits_control(ld_48_io_enable_bits_control),
    .io_Out_0_ready(ld_48_io_Out_0_ready),
    .io_Out_0_valid(ld_48_io_Out_0_valid),
    .io_Out_0_bits_data(ld_48_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_48_io_GepAddr_ready),
    .io_GepAddr_valid(ld_48_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_48_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_48_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_48_io_GepAddr_bits_data),
    .io_memReq_ready(ld_48_io_memReq_ready),
    .io_memReq_valid(ld_48_io_memReq_valid),
    .io_memReq_bits_address(ld_48_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_48_io_memReq_bits_taskID),
    .io_memResp_valid(ld_48_io_memResp_valid),
    .io_memResp_data(ld_48_io_memResp_data)
  );
  ComputeNode_22 binaryOp_add4249 ( // @[extracted_function_conv.scala 236:32]
    .clock(binaryOp_add4249_clock),
    .reset(binaryOp_add4249_reset),
    .io_enable_ready(binaryOp_add4249_io_enable_ready),
    .io_enable_valid(binaryOp_add4249_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add4249_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add4249_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add4249_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add4249_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add4249_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add4249_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add4249_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add4249_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add4249_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add4249_io_RightIO_valid)
  );
  GepNode_11 Gep_arrayidx4350 ( // @[extracted_function_conv.scala 239:32]
    .clock(Gep_arrayidx4350_clock),
    .reset(Gep_arrayidx4350_reset),
    .io_enable_ready(Gep_arrayidx4350_io_enable_ready),
    .io_enable_valid(Gep_arrayidx4350_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx4350_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx4350_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx4350_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx4350_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx4350_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx4350_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx4350_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx4350_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx4350_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx4350_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx4350_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx4350_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx4350_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx4350_io_idx_0_bits_data)
  );
  UnTypLoad_6 ld_51 ( // @[extracted_function_conv.scala 242:21]
    .clock(ld_51_clock),
    .reset(ld_51_reset),
    .io_enable_ready(ld_51_io_enable_ready),
    .io_enable_valid(ld_51_io_enable_valid),
    .io_enable_bits_taskID(ld_51_io_enable_bits_taskID),
    .io_enable_bits_control(ld_51_io_enable_bits_control),
    .io_Out_0_ready(ld_51_io_Out_0_ready),
    .io_Out_0_valid(ld_51_io_Out_0_valid),
    .io_Out_0_bits_data(ld_51_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_51_io_GepAddr_ready),
    .io_GepAddr_valid(ld_51_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_51_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_51_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_51_io_GepAddr_bits_data),
    .io_memReq_ready(ld_51_io_memReq_ready),
    .io_memReq_valid(ld_51_io_memReq_valid),
    .io_memReq_bits_address(ld_51_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_51_io_memReq_bits_taskID),
    .io_memResp_valid(ld_51_io_memResp_valid),
    .io_memResp_data(ld_51_io_memResp_data)
  );
  ZextNode_2 sextconv4552 ( // @[extracted_function_conv.scala 245:28]
    .clock(sextconv4552_clock),
    .reset(sextconv4552_reset),
    .io_Input_ready(sextconv4552_io_Input_ready),
    .io_Input_valid(sextconv4552_io_Input_valid),
    .io_Input_bits_data(sextconv4552_io_Input_bits_data),
    .io_enable_ready(sextconv4552_io_enable_ready),
    .io_enable_valid(sextconv4552_io_enable_valid),
    .io_enable_bits_taskID(sextconv4552_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv4552_io_Out_0_ready),
    .io_Out_0_valid(sextconv4552_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv4552_io_Out_0_bits_data)
  );
  ComputeNode_23 binaryOp_mul4653 ( // @[extracted_function_conv.scala 248:32]
    .clock(binaryOp_mul4653_clock),
    .reset(binaryOp_mul4653_reset),
    .io_enable_ready(binaryOp_mul4653_io_enable_ready),
    .io_enable_valid(binaryOp_mul4653_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul4653_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul4653_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul4653_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul4653_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul4653_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul4653_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul4653_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul4653_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul4653_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul4653_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul4653_io_RightIO_bits_data)
  );
  ComputeNode_24 binaryOp_add4754 ( // @[extracted_function_conv.scala 251:32]
    .clock(binaryOp_add4754_clock),
    .reset(binaryOp_add4754_reset),
    .io_enable_ready(binaryOp_add4754_io_enable_ready),
    .io_enable_valid(binaryOp_add4754_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add4754_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add4754_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add4754_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add4754_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add4754_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add4754_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add4754_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add4754_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add4754_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add4754_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add4754_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add4754_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add4754_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add4754_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add4754_io_RightIO_bits_data)
  );
  UnTypStore_2 st_55 ( // @[extracted_function_conv.scala 254:21]
    .clock(st_55_clock),
    .reset(st_55_reset),
    .io_enable_ready(st_55_io_enable_ready),
    .io_enable_valid(st_55_io_enable_valid),
    .io_enable_bits_taskID(st_55_io_enable_bits_taskID),
    .io_enable_bits_control(st_55_io_enable_bits_control),
    .io_GepAddr_ready(st_55_io_GepAddr_ready),
    .io_GepAddr_valid(st_55_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_55_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_55_io_GepAddr_bits_data),
    .io_inData_ready(st_55_io_inData_ready),
    .io_inData_valid(st_55_io_inData_valid),
    .io_inData_bits_taskID(st_55_io_inData_bits_taskID),
    .io_inData_bits_data(st_55_io_inData_bits_data),
    .io_memReq_ready(st_55_io_memReq_ready),
    .io_memReq_valid(st_55_io_memReq_valid),
    .io_memReq_bits_address(st_55_io_memReq_bits_address),
    .io_memReq_bits_data(st_55_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_55_io_memReq_bits_taskID),
    .io_memResp_valid(st_55_io_memResp_valid)
  );
  UnTypLoad_7 ld_56 ( // @[extracted_function_conv.scala 257:21]
    .clock(ld_56_clock),
    .reset(ld_56_reset),
    .io_enable_ready(ld_56_io_enable_ready),
    .io_enable_valid(ld_56_io_enable_valid),
    .io_enable_bits_taskID(ld_56_io_enable_bits_taskID),
    .io_enable_bits_control(ld_56_io_enable_bits_control),
    .io_Out_0_ready(ld_56_io_Out_0_ready),
    .io_Out_0_valid(ld_56_io_Out_0_valid),
    .io_Out_0_bits_data(ld_56_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_56_io_GepAddr_ready),
    .io_GepAddr_valid(ld_56_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_56_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_56_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_56_io_GepAddr_bits_data),
    .io_memReq_ready(ld_56_io_memReq_ready),
    .io_memReq_valid(ld_56_io_memReq_valid),
    .io_memReq_bits_address(ld_56_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_56_io_memReq_bits_taskID),
    .io_memResp_valid(ld_56_io_memResp_valid),
    .io_memResp_data(ld_56_io_memResp_data)
  );
  ComputeNode_25 binaryOp_mul5257 ( // @[extracted_function_conv.scala 260:32]
    .clock(binaryOp_mul5257_clock),
    .reset(binaryOp_mul5257_reset),
    .io_enable_ready(binaryOp_mul5257_io_enable_ready),
    .io_enable_valid(binaryOp_mul5257_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul5257_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul5257_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul5257_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul5257_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul5257_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_mul5257_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_mul5257_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_mul5257_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_mul5257_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul5257_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul5257_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul5257_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul5257_io_RightIO_valid)
  );
  ComputeNode_26 binaryOp_add5358 ( // @[extracted_function_conv.scala 263:32]
    .clock(binaryOp_add5358_clock),
    .reset(binaryOp_add5358_reset),
    .io_enable_ready(binaryOp_add5358_io_enable_ready),
    .io_enable_valid(binaryOp_add5358_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add5358_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add5358_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add5358_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add5358_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add5358_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add5358_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add5358_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add5358_io_Out_1_bits_data),
    .io_Out_2_ready(binaryOp_add5358_io_Out_2_ready),
    .io_Out_2_valid(binaryOp_add5358_io_Out_2_valid),
    .io_Out_2_bits_data(binaryOp_add5358_io_Out_2_bits_data),
    .io_LeftIO_ready(binaryOp_add5358_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add5358_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add5358_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add5358_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add5358_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add5358_io_RightIO_bits_data)
  );
  GepNode_12 Gep_arrayidx5459 ( // @[extracted_function_conv.scala 266:32]
    .clock(Gep_arrayidx5459_clock),
    .reset(Gep_arrayidx5459_reset),
    .io_enable_ready(Gep_arrayidx5459_io_enable_ready),
    .io_enable_valid(Gep_arrayidx5459_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx5459_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx5459_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx5459_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx5459_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx5459_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx5459_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx5459_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx5459_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx5459_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx5459_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx5459_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx5459_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx5459_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx5459_io_idx_0_bits_data)
  );
  UnTypLoad_8 ld_60 ( // @[extracted_function_conv.scala 269:21]
    .clock(ld_60_clock),
    .reset(ld_60_reset),
    .io_enable_ready(ld_60_io_enable_ready),
    .io_enable_valid(ld_60_io_enable_valid),
    .io_enable_bits_taskID(ld_60_io_enable_bits_taskID),
    .io_enable_bits_control(ld_60_io_enable_bits_control),
    .io_Out_0_ready(ld_60_io_Out_0_ready),
    .io_Out_0_valid(ld_60_io_Out_0_valid),
    .io_Out_0_bits_data(ld_60_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_60_io_GepAddr_ready),
    .io_GepAddr_valid(ld_60_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_60_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_60_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_60_io_GepAddr_bits_data),
    .io_memReq_ready(ld_60_io_memReq_ready),
    .io_memReq_valid(ld_60_io_memReq_valid),
    .io_memReq_bits_address(ld_60_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_60_io_memReq_bits_taskID),
    .io_memResp_valid(ld_60_io_memResp_valid),
    .io_memResp_data(ld_60_io_memResp_data)
  );
  ZextNode_3 sextconv5661 ( // @[extracted_function_conv.scala 272:28]
    .clock(sextconv5661_clock),
    .reset(sextconv5661_reset),
    .io_Input_ready(sextconv5661_io_Input_ready),
    .io_Input_valid(sextconv5661_io_Input_valid),
    .io_Input_bits_data(sextconv5661_io_Input_bits_data),
    .io_enable_ready(sextconv5661_io_enable_ready),
    .io_enable_valid(sextconv5661_io_enable_valid),
    .io_enable_bits_taskID(sextconv5661_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv5661_io_Out_0_ready),
    .io_Out_0_valid(sextconv5661_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv5661_io_Out_0_bits_data)
  );
  ComputeNode_27 binaryOp_mul5762 ( // @[extracted_function_conv.scala 275:32]
    .clock(binaryOp_mul5762_clock),
    .reset(binaryOp_mul5762_reset),
    .io_enable_ready(binaryOp_mul5762_io_enable_ready),
    .io_enable_valid(binaryOp_mul5762_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul5762_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul5762_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul5762_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul5762_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul5762_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul5762_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul5762_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul5762_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul5762_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul5762_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul5762_io_RightIO_bits_data)
  );
  ComputeNode_28 binaryOp_add5863 ( // @[extracted_function_conv.scala 278:32]
    .clock(binaryOp_add5863_clock),
    .reset(binaryOp_add5863_reset),
    .io_enable_ready(binaryOp_add5863_io_enable_ready),
    .io_enable_valid(binaryOp_add5863_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add5863_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add5863_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add5863_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add5863_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add5863_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add5863_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add5863_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add5863_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add5863_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add5863_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add5863_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add5863_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add5863_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add5863_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add5863_io_RightIO_bits_data)
  );
  UnTypStore_3 st_64 ( // @[extracted_function_conv.scala 281:21]
    .clock(st_64_clock),
    .reset(st_64_reset),
    .io_enable_ready(st_64_io_enable_ready),
    .io_enable_valid(st_64_io_enable_valid),
    .io_enable_bits_taskID(st_64_io_enable_bits_taskID),
    .io_enable_bits_control(st_64_io_enable_bits_control),
    .io_GepAddr_ready(st_64_io_GepAddr_ready),
    .io_GepAddr_valid(st_64_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_64_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_64_io_GepAddr_bits_data),
    .io_inData_ready(st_64_io_inData_ready),
    .io_inData_valid(st_64_io_inData_valid),
    .io_inData_bits_taskID(st_64_io_inData_bits_taskID),
    .io_inData_bits_data(st_64_io_inData_bits_data),
    .io_memReq_ready(st_64_io_memReq_ready),
    .io_memReq_valid(st_64_io_memReq_valid),
    .io_memReq_bits_address(st_64_io_memReq_bits_address),
    .io_memReq_bits_data(st_64_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_64_io_memReq_bits_taskID),
    .io_memResp_valid(st_64_io_memResp_valid)
  );
  UnTypLoad_9 ld_65 ( // @[extracted_function_conv.scala 284:21]
    .clock(ld_65_clock),
    .reset(ld_65_reset),
    .io_enable_ready(ld_65_io_enable_ready),
    .io_enable_valid(ld_65_io_enable_valid),
    .io_enable_bits_taskID(ld_65_io_enable_bits_taskID),
    .io_enable_bits_control(ld_65_io_enable_bits_control),
    .io_Out_0_ready(ld_65_io_Out_0_ready),
    .io_Out_0_valid(ld_65_io_Out_0_valid),
    .io_Out_0_bits_data(ld_65_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_65_io_GepAddr_ready),
    .io_GepAddr_valid(ld_65_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_65_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_65_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_65_io_GepAddr_bits_data),
    .io_memReq_ready(ld_65_io_memReq_ready),
    .io_memReq_valid(ld_65_io_memReq_valid),
    .io_memReq_bits_address(ld_65_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_65_io_memReq_bits_taskID),
    .io_memResp_valid(ld_65_io_memResp_valid),
    .io_memResp_data(ld_65_io_memResp_data)
  );
  ComputeNode_29 binaryOp_add6566 ( // @[extracted_function_conv.scala 287:32]
    .clock(binaryOp_add6566_clock),
    .reset(binaryOp_add6566_reset),
    .io_enable_ready(binaryOp_add6566_io_enable_ready),
    .io_enable_valid(binaryOp_add6566_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add6566_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add6566_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add6566_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add6566_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add6566_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add6566_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add6566_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add6566_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add6566_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add6566_io_RightIO_valid)
  );
  GepNode_13 Gep_arrayidx6667 ( // @[extracted_function_conv.scala 290:32]
    .clock(Gep_arrayidx6667_clock),
    .reset(Gep_arrayidx6667_reset),
    .io_enable_ready(Gep_arrayidx6667_io_enable_ready),
    .io_enable_valid(Gep_arrayidx6667_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx6667_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx6667_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx6667_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx6667_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx6667_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx6667_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx6667_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx6667_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx6667_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx6667_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx6667_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx6667_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx6667_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx6667_io_idx_0_bits_data)
  );
  UnTypLoad_10 ld_68 ( // @[extracted_function_conv.scala 293:21]
    .clock(ld_68_clock),
    .reset(ld_68_reset),
    .io_enable_ready(ld_68_io_enable_ready),
    .io_enable_valid(ld_68_io_enable_valid),
    .io_enable_bits_taskID(ld_68_io_enable_bits_taskID),
    .io_enable_bits_control(ld_68_io_enable_bits_control),
    .io_Out_0_ready(ld_68_io_Out_0_ready),
    .io_Out_0_valid(ld_68_io_Out_0_valid),
    .io_Out_0_bits_data(ld_68_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_68_io_GepAddr_ready),
    .io_GepAddr_valid(ld_68_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_68_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_68_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_68_io_GepAddr_bits_data),
    .io_memReq_ready(ld_68_io_memReq_ready),
    .io_memReq_valid(ld_68_io_memReq_valid),
    .io_memReq_bits_address(ld_68_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_68_io_memReq_bits_taskID),
    .io_memResp_valid(ld_68_io_memResp_valid),
    .io_memResp_data(ld_68_io_memResp_data)
  );
  ZextNode_4 sextconv6869 ( // @[extracted_function_conv.scala 296:28]
    .clock(sextconv6869_clock),
    .reset(sextconv6869_reset),
    .io_Input_ready(sextconv6869_io_Input_ready),
    .io_Input_valid(sextconv6869_io_Input_valid),
    .io_Input_bits_data(sextconv6869_io_Input_bits_data),
    .io_enable_ready(sextconv6869_io_enable_ready),
    .io_enable_valid(sextconv6869_io_enable_valid),
    .io_enable_bits_taskID(sextconv6869_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv6869_io_Out_0_ready),
    .io_Out_0_valid(sextconv6869_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv6869_io_Out_0_bits_data)
  );
  ComputeNode_30 binaryOp_mul6970 ( // @[extracted_function_conv.scala 299:32]
    .clock(binaryOp_mul6970_clock),
    .reset(binaryOp_mul6970_reset),
    .io_enable_ready(binaryOp_mul6970_io_enable_ready),
    .io_enable_valid(binaryOp_mul6970_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul6970_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul6970_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul6970_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul6970_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul6970_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul6970_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul6970_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul6970_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul6970_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul6970_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul6970_io_RightIO_bits_data)
  );
  ComputeNode_31 binaryOp_add7071 ( // @[extracted_function_conv.scala 302:32]
    .clock(binaryOp_add7071_clock),
    .reset(binaryOp_add7071_reset),
    .io_enable_ready(binaryOp_add7071_io_enable_ready),
    .io_enable_valid(binaryOp_add7071_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add7071_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add7071_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add7071_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add7071_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add7071_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add7071_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add7071_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add7071_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add7071_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add7071_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add7071_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add7071_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add7071_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add7071_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add7071_io_RightIO_bits_data)
  );
  UnTypStore_4 st_72 ( // @[extracted_function_conv.scala 305:21]
    .clock(st_72_clock),
    .reset(st_72_reset),
    .io_enable_ready(st_72_io_enable_ready),
    .io_enable_valid(st_72_io_enable_valid),
    .io_enable_bits_taskID(st_72_io_enable_bits_taskID),
    .io_enable_bits_control(st_72_io_enable_bits_control),
    .io_GepAddr_ready(st_72_io_GepAddr_ready),
    .io_GepAddr_valid(st_72_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_72_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_72_io_GepAddr_bits_data),
    .io_inData_ready(st_72_io_inData_ready),
    .io_inData_valid(st_72_io_inData_valid),
    .io_inData_bits_taskID(st_72_io_inData_bits_taskID),
    .io_inData_bits_data(st_72_io_inData_bits_data),
    .io_memReq_ready(st_72_io_memReq_ready),
    .io_memReq_valid(st_72_io_memReq_valid),
    .io_memReq_bits_address(st_72_io_memReq_bits_address),
    .io_memReq_bits_data(st_72_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_72_io_memReq_bits_taskID),
    .io_memResp_valid(st_72_io_memResp_valid)
  );
  UnTypLoad_11 ld_73 ( // @[extracted_function_conv.scala 308:21]
    .clock(ld_73_clock),
    .reset(ld_73_reset),
    .io_enable_ready(ld_73_io_enable_ready),
    .io_enable_valid(ld_73_io_enable_valid),
    .io_enable_bits_taskID(ld_73_io_enable_bits_taskID),
    .io_enable_bits_control(ld_73_io_enable_bits_control),
    .io_Out_0_ready(ld_73_io_Out_0_ready),
    .io_Out_0_valid(ld_73_io_Out_0_valid),
    .io_Out_0_bits_data(ld_73_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_73_io_GepAddr_ready),
    .io_GepAddr_valid(ld_73_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_73_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_73_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_73_io_GepAddr_bits_data),
    .io_memReq_ready(ld_73_io_memReq_ready),
    .io_memReq_valid(ld_73_io_memReq_valid),
    .io_memReq_bits_address(ld_73_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_73_io_memReq_bits_taskID),
    .io_memResp_valid(ld_73_io_memResp_valid),
    .io_memResp_data(ld_73_io_memResp_data)
  );
  ComputeNode_32 binaryOp_add7774 ( // @[extracted_function_conv.scala 311:32]
    .clock(binaryOp_add7774_clock),
    .reset(binaryOp_add7774_reset),
    .io_enable_ready(binaryOp_add7774_io_enable_ready),
    .io_enable_valid(binaryOp_add7774_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add7774_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add7774_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add7774_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add7774_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add7774_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add7774_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add7774_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add7774_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add7774_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add7774_io_RightIO_valid)
  );
  GepNode_14 Gep_arrayidx7875 ( // @[extracted_function_conv.scala 314:32]
    .clock(Gep_arrayidx7875_clock),
    .reset(Gep_arrayidx7875_reset),
    .io_enable_ready(Gep_arrayidx7875_io_enable_ready),
    .io_enable_valid(Gep_arrayidx7875_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx7875_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx7875_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx7875_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx7875_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx7875_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx7875_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx7875_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx7875_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx7875_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx7875_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx7875_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx7875_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx7875_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx7875_io_idx_0_bits_data)
  );
  UnTypLoad_12 ld_76 ( // @[extracted_function_conv.scala 317:21]
    .clock(ld_76_clock),
    .reset(ld_76_reset),
    .io_enable_ready(ld_76_io_enable_ready),
    .io_enable_valid(ld_76_io_enable_valid),
    .io_enable_bits_taskID(ld_76_io_enable_bits_taskID),
    .io_enable_bits_control(ld_76_io_enable_bits_control),
    .io_Out_0_ready(ld_76_io_Out_0_ready),
    .io_Out_0_valid(ld_76_io_Out_0_valid),
    .io_Out_0_bits_data(ld_76_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_76_io_GepAddr_ready),
    .io_GepAddr_valid(ld_76_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_76_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_76_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_76_io_GepAddr_bits_data),
    .io_memReq_ready(ld_76_io_memReq_ready),
    .io_memReq_valid(ld_76_io_memReq_valid),
    .io_memReq_bits_address(ld_76_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_76_io_memReq_bits_taskID),
    .io_memResp_valid(ld_76_io_memResp_valid),
    .io_memResp_data(ld_76_io_memResp_data)
  );
  ZextNode_5 sextconv8077 ( // @[extracted_function_conv.scala 320:28]
    .clock(sextconv8077_clock),
    .reset(sextconv8077_reset),
    .io_Input_ready(sextconv8077_io_Input_ready),
    .io_Input_valid(sextconv8077_io_Input_valid),
    .io_Input_bits_data(sextconv8077_io_Input_bits_data),
    .io_enable_ready(sextconv8077_io_enable_ready),
    .io_enable_valid(sextconv8077_io_enable_valid),
    .io_enable_bits_taskID(sextconv8077_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv8077_io_Out_0_ready),
    .io_Out_0_valid(sextconv8077_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv8077_io_Out_0_bits_data)
  );
  ComputeNode_33 binaryOp_mul8178 ( // @[extracted_function_conv.scala 323:32]
    .clock(binaryOp_mul8178_clock),
    .reset(binaryOp_mul8178_reset),
    .io_enable_ready(binaryOp_mul8178_io_enable_ready),
    .io_enable_valid(binaryOp_mul8178_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul8178_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul8178_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul8178_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul8178_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul8178_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul8178_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul8178_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul8178_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul8178_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul8178_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul8178_io_RightIO_bits_data)
  );
  ComputeNode_34 binaryOp_add8279 ( // @[extracted_function_conv.scala 326:32]
    .clock(binaryOp_add8279_clock),
    .reset(binaryOp_add8279_reset),
    .io_enable_ready(binaryOp_add8279_io_enable_ready),
    .io_enable_valid(binaryOp_add8279_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add8279_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add8279_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add8279_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add8279_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add8279_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add8279_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add8279_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add8279_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add8279_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add8279_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add8279_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add8279_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add8279_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add8279_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add8279_io_RightIO_bits_data)
  );
  UnTypStore_5 st_80 ( // @[extracted_function_conv.scala 329:21]
    .clock(st_80_clock),
    .reset(st_80_reset),
    .io_enable_ready(st_80_io_enable_ready),
    .io_enable_valid(st_80_io_enable_valid),
    .io_enable_bits_taskID(st_80_io_enable_bits_taskID),
    .io_enable_bits_control(st_80_io_enable_bits_control),
    .io_GepAddr_ready(st_80_io_GepAddr_ready),
    .io_GepAddr_valid(st_80_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_80_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_80_io_GepAddr_bits_data),
    .io_inData_ready(st_80_io_inData_ready),
    .io_inData_valid(st_80_io_inData_valid),
    .io_inData_bits_taskID(st_80_io_inData_bits_taskID),
    .io_inData_bits_data(st_80_io_inData_bits_data),
    .io_memReq_ready(st_80_io_memReq_ready),
    .io_memReq_valid(st_80_io_memReq_valid),
    .io_memReq_bits_address(st_80_io_memReq_bits_address),
    .io_memReq_bits_data(st_80_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_80_io_memReq_bits_taskID),
    .io_memResp_valid(st_80_io_memResp_valid)
  );
  UnTypLoad_13 ld_81 ( // @[extracted_function_conv.scala 332:21]
    .clock(ld_81_clock),
    .reset(ld_81_reset),
    .io_enable_ready(ld_81_io_enable_ready),
    .io_enable_valid(ld_81_io_enable_valid),
    .io_enable_bits_taskID(ld_81_io_enable_bits_taskID),
    .io_enable_bits_control(ld_81_io_enable_bits_control),
    .io_Out_0_ready(ld_81_io_Out_0_ready),
    .io_Out_0_valid(ld_81_io_Out_0_valid),
    .io_Out_0_bits_data(ld_81_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_81_io_GepAddr_ready),
    .io_GepAddr_valid(ld_81_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_81_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_81_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_81_io_GepAddr_bits_data),
    .io_memReq_ready(ld_81_io_memReq_ready),
    .io_memReq_valid(ld_81_io_memReq_valid),
    .io_memReq_bits_address(ld_81_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_81_io_memReq_bits_taskID),
    .io_memResp_valid(ld_81_io_memResp_valid),
    .io_memResp_data(ld_81_io_memResp_data)
  );
  ComputeNode_35 binaryOp_add8882 ( // @[extracted_function_conv.scala 335:32]
    .clock(binaryOp_add8882_clock),
    .reset(binaryOp_add8882_reset),
    .io_enable_ready(binaryOp_add8882_io_enable_ready),
    .io_enable_valid(binaryOp_add8882_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add8882_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add8882_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add8882_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add8882_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add8882_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add8882_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add8882_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add8882_io_Out_1_bits_data),
    .io_Out_2_ready(binaryOp_add8882_io_Out_2_ready),
    .io_Out_2_valid(binaryOp_add8882_io_Out_2_valid),
    .io_Out_2_bits_data(binaryOp_add8882_io_Out_2_bits_data),
    .io_LeftIO_ready(binaryOp_add8882_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add8882_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add8882_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add8882_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add8882_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add8882_io_RightIO_bits_data)
  );
  GepNode_15 Gep_arrayidx8983 ( // @[extracted_function_conv.scala 338:32]
    .clock(Gep_arrayidx8983_clock),
    .reset(Gep_arrayidx8983_reset),
    .io_enable_ready(Gep_arrayidx8983_io_enable_ready),
    .io_enable_valid(Gep_arrayidx8983_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx8983_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx8983_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx8983_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx8983_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx8983_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx8983_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx8983_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx8983_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx8983_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx8983_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx8983_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx8983_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx8983_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx8983_io_idx_0_bits_data)
  );
  UnTypLoad_14 ld_84 ( // @[extracted_function_conv.scala 341:21]
    .clock(ld_84_clock),
    .reset(ld_84_reset),
    .io_enable_ready(ld_84_io_enable_ready),
    .io_enable_valid(ld_84_io_enable_valid),
    .io_enable_bits_taskID(ld_84_io_enable_bits_taskID),
    .io_enable_bits_control(ld_84_io_enable_bits_control),
    .io_Out_0_ready(ld_84_io_Out_0_ready),
    .io_Out_0_valid(ld_84_io_Out_0_valid),
    .io_Out_0_bits_data(ld_84_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_84_io_GepAddr_ready),
    .io_GepAddr_valid(ld_84_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_84_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_84_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_84_io_GepAddr_bits_data),
    .io_memReq_ready(ld_84_io_memReq_ready),
    .io_memReq_valid(ld_84_io_memReq_valid),
    .io_memReq_bits_address(ld_84_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_84_io_memReq_bits_taskID),
    .io_memResp_valid(ld_84_io_memResp_valid),
    .io_memResp_data(ld_84_io_memResp_data)
  );
  ZextNode_6 sextconv9185 ( // @[extracted_function_conv.scala 344:28]
    .clock(sextconv9185_clock),
    .reset(sextconv9185_reset),
    .io_Input_ready(sextconv9185_io_Input_ready),
    .io_Input_valid(sextconv9185_io_Input_valid),
    .io_Input_bits_data(sextconv9185_io_Input_bits_data),
    .io_enable_ready(sextconv9185_io_enable_ready),
    .io_enable_valid(sextconv9185_io_enable_valid),
    .io_enable_bits_taskID(sextconv9185_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv9185_io_Out_0_ready),
    .io_Out_0_valid(sextconv9185_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv9185_io_Out_0_bits_data)
  );
  ComputeNode_36 binaryOp_mul9286 ( // @[extracted_function_conv.scala 347:32]
    .clock(binaryOp_mul9286_clock),
    .reset(binaryOp_mul9286_reset),
    .io_enable_ready(binaryOp_mul9286_io_enable_ready),
    .io_enable_valid(binaryOp_mul9286_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul9286_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul9286_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul9286_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul9286_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul9286_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul9286_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul9286_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul9286_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul9286_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul9286_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul9286_io_RightIO_bits_data)
  );
  ComputeNode_37 binaryOp_add9387 ( // @[extracted_function_conv.scala 350:32]
    .clock(binaryOp_add9387_clock),
    .reset(binaryOp_add9387_reset),
    .io_enable_ready(binaryOp_add9387_io_enable_ready),
    .io_enable_valid(binaryOp_add9387_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add9387_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add9387_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add9387_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add9387_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add9387_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add9387_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add9387_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add9387_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add9387_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add9387_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add9387_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add9387_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add9387_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add9387_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add9387_io_RightIO_bits_data)
  );
  UnTypStore_6 st_88 ( // @[extracted_function_conv.scala 353:21]
    .clock(st_88_clock),
    .reset(st_88_reset),
    .io_enable_ready(st_88_io_enable_ready),
    .io_enable_valid(st_88_io_enable_valid),
    .io_enable_bits_taskID(st_88_io_enable_bits_taskID),
    .io_enable_bits_control(st_88_io_enable_bits_control),
    .io_GepAddr_ready(st_88_io_GepAddr_ready),
    .io_GepAddr_valid(st_88_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_88_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_88_io_GepAddr_bits_data),
    .io_inData_ready(st_88_io_inData_ready),
    .io_inData_valid(st_88_io_inData_valid),
    .io_inData_bits_taskID(st_88_io_inData_bits_taskID),
    .io_inData_bits_data(st_88_io_inData_bits_data),
    .io_memReq_ready(st_88_io_memReq_ready),
    .io_memReq_valid(st_88_io_memReq_valid),
    .io_memReq_bits_address(st_88_io_memReq_bits_address),
    .io_memReq_bits_data(st_88_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_88_io_memReq_bits_taskID),
    .io_memResp_valid(st_88_io_memResp_valid)
  );
  UnTypLoad_15 ld_89 ( // @[extracted_function_conv.scala 356:21]
    .clock(ld_89_clock),
    .reset(ld_89_reset),
    .io_enable_ready(ld_89_io_enable_ready),
    .io_enable_valid(ld_89_io_enable_valid),
    .io_enable_bits_taskID(ld_89_io_enable_bits_taskID),
    .io_enable_bits_control(ld_89_io_enable_bits_control),
    .io_Out_0_ready(ld_89_io_Out_0_ready),
    .io_Out_0_valid(ld_89_io_Out_0_valid),
    .io_Out_0_bits_data(ld_89_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_89_io_GepAddr_ready),
    .io_GepAddr_valid(ld_89_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_89_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_89_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_89_io_GepAddr_bits_data),
    .io_memReq_ready(ld_89_io_memReq_ready),
    .io_memReq_valid(ld_89_io_memReq_valid),
    .io_memReq_bits_address(ld_89_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_89_io_memReq_bits_taskID),
    .io_memResp_valid(ld_89_io_memResp_valid),
    .io_memResp_data(ld_89_io_memResp_data)
  );
  ComputeNode_38 binaryOp_add10090 ( // @[extracted_function_conv.scala 359:33]
    .clock(binaryOp_add10090_clock),
    .reset(binaryOp_add10090_reset),
    .io_enable_ready(binaryOp_add10090_io_enable_ready),
    .io_enable_valid(binaryOp_add10090_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add10090_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add10090_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add10090_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add10090_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add10090_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add10090_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add10090_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add10090_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add10090_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add10090_io_RightIO_valid)
  );
  GepNode_16 Gep_arrayidx10191 ( // @[extracted_function_conv.scala 362:33]
    .clock(Gep_arrayidx10191_clock),
    .reset(Gep_arrayidx10191_reset),
    .io_enable_ready(Gep_arrayidx10191_io_enable_ready),
    .io_enable_valid(Gep_arrayidx10191_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx10191_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx10191_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx10191_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx10191_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx10191_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx10191_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx10191_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx10191_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx10191_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx10191_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx10191_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx10191_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx10191_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx10191_io_idx_0_bits_data)
  );
  UnTypLoad_16 ld_92 ( // @[extracted_function_conv.scala 365:21]
    .clock(ld_92_clock),
    .reset(ld_92_reset),
    .io_enable_ready(ld_92_io_enable_ready),
    .io_enable_valid(ld_92_io_enable_valid),
    .io_enable_bits_taskID(ld_92_io_enable_bits_taskID),
    .io_enable_bits_control(ld_92_io_enable_bits_control),
    .io_Out_0_ready(ld_92_io_Out_0_ready),
    .io_Out_0_valid(ld_92_io_Out_0_valid),
    .io_Out_0_bits_data(ld_92_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_92_io_GepAddr_ready),
    .io_GepAddr_valid(ld_92_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_92_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_92_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_92_io_GepAddr_bits_data),
    .io_memReq_ready(ld_92_io_memReq_ready),
    .io_memReq_valid(ld_92_io_memReq_valid),
    .io_memReq_bits_address(ld_92_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_92_io_memReq_bits_taskID),
    .io_memResp_valid(ld_92_io_memResp_valid),
    .io_memResp_data(ld_92_io_memResp_data)
  );
  ZextNode_7 sextconv10393 ( // @[extracted_function_conv.scala 368:29]
    .clock(sextconv10393_clock),
    .reset(sextconv10393_reset),
    .io_Input_ready(sextconv10393_io_Input_ready),
    .io_Input_valid(sextconv10393_io_Input_valid),
    .io_Input_bits_data(sextconv10393_io_Input_bits_data),
    .io_enable_ready(sextconv10393_io_enable_ready),
    .io_enable_valid(sextconv10393_io_enable_valid),
    .io_enable_bits_taskID(sextconv10393_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv10393_io_Out_0_ready),
    .io_Out_0_valid(sextconv10393_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv10393_io_Out_0_bits_data)
  );
  ComputeNode_39 binaryOp_mul10494 ( // @[extracted_function_conv.scala 371:33]
    .clock(binaryOp_mul10494_clock),
    .reset(binaryOp_mul10494_reset),
    .io_enable_ready(binaryOp_mul10494_io_enable_ready),
    .io_enable_valid(binaryOp_mul10494_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul10494_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul10494_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul10494_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul10494_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul10494_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul10494_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul10494_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul10494_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul10494_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul10494_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul10494_io_RightIO_bits_data)
  );
  ComputeNode_40 binaryOp_add10595 ( // @[extracted_function_conv.scala 374:33]
    .clock(binaryOp_add10595_clock),
    .reset(binaryOp_add10595_reset),
    .io_enable_ready(binaryOp_add10595_io_enable_ready),
    .io_enable_valid(binaryOp_add10595_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add10595_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add10595_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add10595_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add10595_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add10595_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add10595_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_add10595_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_add10595_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_add10595_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_add10595_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add10595_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add10595_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add10595_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add10595_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add10595_io_RightIO_bits_data)
  );
  UnTypStore_7 st_96 ( // @[extracted_function_conv.scala 377:21]
    .clock(st_96_clock),
    .reset(st_96_reset),
    .io_enable_ready(st_96_io_enable_ready),
    .io_enable_valid(st_96_io_enable_valid),
    .io_enable_bits_taskID(st_96_io_enable_bits_taskID),
    .io_enable_bits_control(st_96_io_enable_bits_control),
    .io_GepAddr_ready(st_96_io_GepAddr_ready),
    .io_GepAddr_valid(st_96_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_96_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_96_io_GepAddr_bits_data),
    .io_inData_ready(st_96_io_inData_ready),
    .io_inData_valid(st_96_io_inData_valid),
    .io_inData_bits_taskID(st_96_io_inData_bits_taskID),
    .io_inData_bits_data(st_96_io_inData_bits_data),
    .io_memReq_ready(st_96_io_memReq_ready),
    .io_memReq_valid(st_96_io_memReq_valid),
    .io_memReq_bits_address(st_96_io_memReq_bits_address),
    .io_memReq_bits_data(st_96_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_96_io_memReq_bits_taskID),
    .io_memResp_valid(st_96_io_memResp_valid)
  );
  UnTypLoad_17 ld_97 ( // @[extracted_function_conv.scala 380:21]
    .clock(ld_97_clock),
    .reset(ld_97_reset),
    .io_enable_ready(ld_97_io_enable_ready),
    .io_enable_valid(ld_97_io_enable_valid),
    .io_enable_bits_taskID(ld_97_io_enable_bits_taskID),
    .io_enable_bits_control(ld_97_io_enable_bits_control),
    .io_Out_0_ready(ld_97_io_Out_0_ready),
    .io_Out_0_valid(ld_97_io_Out_0_valid),
    .io_Out_0_bits_data(ld_97_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_97_io_GepAddr_ready),
    .io_GepAddr_valid(ld_97_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_97_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_97_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_97_io_GepAddr_bits_data),
    .io_memReq_ready(ld_97_io_memReq_ready),
    .io_memReq_valid(ld_97_io_memReq_valid),
    .io_memReq_bits_address(ld_97_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_97_io_memReq_bits_taskID),
    .io_memResp_valid(ld_97_io_memResp_valid),
    .io_memResp_data(ld_97_io_memResp_data)
  );
  ComputeNode_41 binaryOp_add11298 ( // @[extracted_function_conv.scala 383:33]
    .clock(binaryOp_add11298_clock),
    .reset(binaryOp_add11298_reset),
    .io_enable_ready(binaryOp_add11298_io_enable_ready),
    .io_enable_valid(binaryOp_add11298_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add11298_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add11298_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add11298_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add11298_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_add11298_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add11298_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add11298_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add11298_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add11298_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add11298_io_RightIO_valid)
  );
  GepNode_17 Gep_arrayidx11399 ( // @[extracted_function_conv.scala 386:33]
    .clock(Gep_arrayidx11399_clock),
    .reset(Gep_arrayidx11399_reset),
    .io_enable_ready(Gep_arrayidx11399_io_enable_ready),
    .io_enable_valid(Gep_arrayidx11399_io_enable_valid),
    .io_enable_bits_taskID(Gep_arrayidx11399_io_enable_bits_taskID),
    .io_enable_bits_control(Gep_arrayidx11399_io_enable_bits_control),
    .io_Out_0_ready(Gep_arrayidx11399_io_Out_0_ready),
    .io_Out_0_valid(Gep_arrayidx11399_io_Out_0_valid),
    .io_Out_0_bits_predicate(Gep_arrayidx11399_io_Out_0_bits_predicate),
    .io_Out_0_bits_taskID(Gep_arrayidx11399_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(Gep_arrayidx11399_io_Out_0_bits_data),
    .io_baseAddress_ready(Gep_arrayidx11399_io_baseAddress_ready),
    .io_baseAddress_valid(Gep_arrayidx11399_io_baseAddress_valid),
    .io_baseAddress_bits_taskID(Gep_arrayidx11399_io_baseAddress_bits_taskID),
    .io_baseAddress_bits_data(Gep_arrayidx11399_io_baseAddress_bits_data),
    .io_idx_0_ready(Gep_arrayidx11399_io_idx_0_ready),
    .io_idx_0_valid(Gep_arrayidx11399_io_idx_0_valid),
    .io_idx_0_bits_data(Gep_arrayidx11399_io_idx_0_bits_data)
  );
  UnTypLoad_18 ld_100 ( // @[extracted_function_conv.scala 389:22]
    .clock(ld_100_clock),
    .reset(ld_100_reset),
    .io_enable_ready(ld_100_io_enable_ready),
    .io_enable_valid(ld_100_io_enable_valid),
    .io_enable_bits_taskID(ld_100_io_enable_bits_taskID),
    .io_enable_bits_control(ld_100_io_enable_bits_control),
    .io_Out_0_ready(ld_100_io_Out_0_ready),
    .io_Out_0_valid(ld_100_io_Out_0_valid),
    .io_Out_0_bits_data(ld_100_io_Out_0_bits_data),
    .io_GepAddr_ready(ld_100_io_GepAddr_ready),
    .io_GepAddr_valid(ld_100_io_GepAddr_valid),
    .io_GepAddr_bits_predicate(ld_100_io_GepAddr_bits_predicate),
    .io_GepAddr_bits_taskID(ld_100_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(ld_100_io_GepAddr_bits_data),
    .io_memReq_ready(ld_100_io_memReq_ready),
    .io_memReq_valid(ld_100_io_memReq_valid),
    .io_memReq_bits_address(ld_100_io_memReq_bits_address),
    .io_memReq_bits_taskID(ld_100_io_memReq_bits_taskID),
    .io_memResp_valid(ld_100_io_memResp_valid),
    .io_memResp_data(ld_100_io_memResp_data)
  );
  ZextNode_8 sextconv115101 ( // @[extracted_function_conv.scala 392:30]
    .clock(sextconv115101_clock),
    .reset(sextconv115101_reset),
    .io_Input_ready(sextconv115101_io_Input_ready),
    .io_Input_valid(sextconv115101_io_Input_valid),
    .io_Input_bits_data(sextconv115101_io_Input_bits_data),
    .io_enable_ready(sextconv115101_io_enable_ready),
    .io_enable_valid(sextconv115101_io_enable_valid),
    .io_enable_bits_taskID(sextconv115101_io_enable_bits_taskID),
    .io_Out_0_ready(sextconv115101_io_Out_0_ready),
    .io_Out_0_valid(sextconv115101_io_Out_0_valid),
    .io_Out_0_bits_data(sextconv115101_io_Out_0_bits_data)
  );
  ComputeNode_42 binaryOp_mul116102 ( // @[extracted_function_conv.scala 395:34]
    .clock(binaryOp_mul116102_clock),
    .reset(binaryOp_mul116102_reset),
    .io_enable_ready(binaryOp_mul116102_io_enable_ready),
    .io_enable_valid(binaryOp_mul116102_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_mul116102_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_mul116102_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_mul116102_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_mul116102_io_Out_0_valid),
    .io_Out_0_bits_data(binaryOp_mul116102_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_mul116102_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_mul116102_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_mul116102_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_mul116102_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_mul116102_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_mul116102_io_RightIO_bits_data)
  );
  ComputeNode_43 binaryOp_add117103 ( // @[extracted_function_conv.scala 398:34]
    .clock(binaryOp_add117103_clock),
    .reset(binaryOp_add117103_reset),
    .io_enable_ready(binaryOp_add117103_io_enable_ready),
    .io_enable_valid(binaryOp_add117103_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_add117103_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_add117103_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_add117103_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_add117103_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_add117103_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_add117103_io_Out_0_bits_data),
    .io_LeftIO_ready(binaryOp_add117103_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_add117103_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_add117103_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_add117103_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_add117103_io_RightIO_valid),
    .io_RightIO_bits_data(binaryOp_add117103_io_RightIO_bits_data)
  );
  UnTypStore_8 st_104 ( // @[extracted_function_conv.scala 401:22]
    .clock(st_104_clock),
    .reset(st_104_reset),
    .io_enable_ready(st_104_io_enable_ready),
    .io_enable_valid(st_104_io_enable_valid),
    .io_enable_bits_taskID(st_104_io_enable_bits_taskID),
    .io_enable_bits_control(st_104_io_enable_bits_control),
    .io_GepAddr_ready(st_104_io_GepAddr_ready),
    .io_GepAddr_valid(st_104_io_GepAddr_valid),
    .io_GepAddr_bits_taskID(st_104_io_GepAddr_bits_taskID),
    .io_GepAddr_bits_data(st_104_io_GepAddr_bits_data),
    .io_inData_ready(st_104_io_inData_ready),
    .io_inData_valid(st_104_io_inData_valid),
    .io_inData_bits_taskID(st_104_io_inData_bits_taskID),
    .io_inData_bits_data(st_104_io_inData_bits_data),
    .io_memReq_ready(st_104_io_memReq_ready),
    .io_memReq_valid(st_104_io_memReq_valid),
    .io_memReq_bits_address(st_104_io_memReq_bits_address),
    .io_memReq_bits_data(st_104_io_memReq_bits_data),
    .io_memReq_bits_taskID(st_104_io_memReq_bits_taskID),
    .io_memResp_valid(st_104_io_memResp_valid)
  );
  ComputeNode_44 binaryOp_inc105 ( // @[extracted_function_conv.scala 404:31]
    .clock(binaryOp_inc105_clock),
    .reset(binaryOp_inc105_reset),
    .io_enable_ready(binaryOp_inc105_io_enable_ready),
    .io_enable_valid(binaryOp_inc105_io_enable_valid),
    .io_enable_bits_taskID(binaryOp_inc105_io_enable_bits_taskID),
    .io_enable_bits_control(binaryOp_inc105_io_enable_bits_control),
    .io_Out_0_ready(binaryOp_inc105_io_Out_0_ready),
    .io_Out_0_valid(binaryOp_inc105_io_Out_0_valid),
    .io_Out_0_bits_taskID(binaryOp_inc105_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(binaryOp_inc105_io_Out_0_bits_data),
    .io_Out_1_ready(binaryOp_inc105_io_Out_1_ready),
    .io_Out_1_valid(binaryOp_inc105_io_Out_1_valid),
    .io_Out_1_bits_data(binaryOp_inc105_io_Out_1_bits_data),
    .io_LeftIO_ready(binaryOp_inc105_io_LeftIO_ready),
    .io_LeftIO_valid(binaryOp_inc105_io_LeftIO_valid),
    .io_LeftIO_bits_data(binaryOp_inc105_io_LeftIO_bits_data),
    .io_RightIO_ready(binaryOp_inc105_io_RightIO_ready),
    .io_RightIO_valid(binaryOp_inc105_io_RightIO_valid)
  );
  ComputeNode_45 icmp_exitcond106 ( // @[extracted_function_conv.scala 407:32]
    .clock(icmp_exitcond106_clock),
    .reset(icmp_exitcond106_reset),
    .io_enable_ready(icmp_exitcond106_io_enable_ready),
    .io_enable_valid(icmp_exitcond106_io_enable_valid),
    .io_enable_bits_taskID(icmp_exitcond106_io_enable_bits_taskID),
    .io_enable_bits_control(icmp_exitcond106_io_enable_bits_control),
    .io_Out_0_ready(icmp_exitcond106_io_Out_0_ready),
    .io_Out_0_valid(icmp_exitcond106_io_Out_0_valid),
    .io_Out_0_bits_taskID(icmp_exitcond106_io_Out_0_bits_taskID),
    .io_Out_0_bits_data(icmp_exitcond106_io_Out_0_bits_data),
    .io_LeftIO_ready(icmp_exitcond106_io_LeftIO_ready),
    .io_LeftIO_valid(icmp_exitcond106_io_LeftIO_valid),
    .io_LeftIO_bits_data(icmp_exitcond106_io_LeftIO_bits_data),
    .io_RightIO_ready(icmp_exitcond106_io_RightIO_ready),
    .io_RightIO_valid(icmp_exitcond106_io_RightIO_valid)
  );
  CBranchNodeVariable_1 br_107 ( // @[extracted_function_conv.scala 410:22]
    .clock(br_107_clock),
    .reset(br_107_reset),
    .io_enable_ready(br_107_io_enable_ready),
    .io_enable_valid(br_107_io_enable_valid),
    .io_enable_bits_taskID(br_107_io_enable_bits_taskID),
    .io_enable_bits_control(br_107_io_enable_bits_control),
    .io_CmpIO_ready(br_107_io_CmpIO_ready),
    .io_CmpIO_valid(br_107_io_CmpIO_valid),
    .io_CmpIO_bits_taskID(br_107_io_CmpIO_bits_taskID),
    .io_CmpIO_bits_data(br_107_io_CmpIO_bits_data),
    .io_TrueOutput_0_ready(br_107_io_TrueOutput_0_ready),
    .io_TrueOutput_0_valid(br_107_io_TrueOutput_0_valid),
    .io_TrueOutput_0_bits_control(br_107_io_TrueOutput_0_bits_control),
    .io_FalseOutput_0_ready(br_107_io_FalseOutput_0_ready),
    .io_FalseOutput_0_valid(br_107_io_FalseOutput_0_valid),
    .io_FalseOutput_0_bits_taskID(br_107_io_FalseOutput_0_bits_taskID),
    .io_FalseOutput_0_bits_control(br_107_io_FalseOutput_0_bits_control)
  );
  ConstFastNode const0 ( // @[extracted_function_conv.scala 419:22]
    .clock(const0_clock),
    .reset(const0_reset),
    .io_enable_ready(const0_io_enable_ready),
    .io_enable_valid(const0_io_enable_valid),
    .io_enable_bits_taskID(const0_io_enable_bits_taskID),
    .io_Out_ready(const0_io_Out_ready),
    .io_Out_valid(const0_io_Out_valid)
  );
  ConstFastNode_1 const1 ( // @[extracted_function_conv.scala 422:22]
    .clock(const1_clock),
    .reset(const1_reset),
    .io_enable_ready(const1_io_enable_ready),
    .io_enable_valid(const1_io_enable_valid),
    .io_enable_bits_taskID(const1_io_enable_bits_taskID),
    .io_Out_ready(const1_io_Out_ready),
    .io_Out_valid(const1_io_Out_valid)
  );
  ConstFastNode_2 const2 ( // @[extracted_function_conv.scala 425:22]
    .clock(const2_clock),
    .reset(const2_reset),
    .io_enable_ready(const2_io_enable_ready),
    .io_enable_valid(const2_io_enable_valid),
    .io_enable_bits_taskID(const2_io_enable_bits_taskID),
    .io_Out_ready(const2_io_Out_ready),
    .io_Out_valid(const2_io_Out_valid)
  );
  ConstFastNode_3 const3 ( // @[extracted_function_conv.scala 428:22]
    .clock(const3_clock),
    .reset(const3_reset),
    .io_enable_ready(const3_io_enable_ready),
    .io_enable_valid(const3_io_enable_valid),
    .io_enable_bits_taskID(const3_io_enable_bits_taskID),
    .io_Out_ready(const3_io_Out_ready),
    .io_Out_valid(const3_io_Out_valid)
  );
  ConstFastNode_4 const4 ( // @[extracted_function_conv.scala 431:22]
    .clock(const4_clock),
    .reset(const4_reset),
    .io_enable_ready(const4_io_enable_ready),
    .io_enable_valid(const4_io_enable_valid),
    .io_enable_bits_taskID(const4_io_enable_bits_taskID),
    .io_Out_ready(const4_io_Out_ready),
    .io_Out_valid(const4_io_Out_valid)
  );
  ConstFastNode_5 const5 ( // @[extracted_function_conv.scala 434:22]
    .clock(const5_clock),
    .reset(const5_reset),
    .io_enable_ready(const5_io_enable_ready),
    .io_enable_valid(const5_io_enable_valid),
    .io_enable_bits_taskID(const5_io_enable_bits_taskID),
    .io_Out_ready(const5_io_Out_ready),
    .io_Out_valid(const5_io_Out_valid)
  );
  ConstFastNode_6 const6 ( // @[extracted_function_conv.scala 437:22]
    .clock(const6_clock),
    .reset(const6_reset),
    .io_enable_ready(const6_io_enable_ready),
    .io_enable_valid(const6_io_enable_valid),
    .io_enable_bits_taskID(const6_io_enable_bits_taskID),
    .io_Out_ready(const6_io_Out_ready),
    .io_Out_valid(const6_io_Out_valid)
  );
  ConstFastNode_7 const7 ( // @[extracted_function_conv.scala 440:22]
    .clock(const7_clock),
    .reset(const7_reset),
    .io_enable_ready(const7_io_enable_ready),
    .io_enable_valid(const7_io_enable_valid),
    .io_enable_bits_taskID(const7_io_enable_bits_taskID),
    .io_Out_ready(const7_io_Out_ready),
    .io_Out_valid(const7_io_Out_valid)
  );
  ConstFastNode_8 const8 ( // @[extracted_function_conv.scala 443:22]
    .clock(const8_clock),
    .reset(const8_reset),
    .io_enable_ready(const8_io_enable_ready),
    .io_enable_valid(const8_io_enable_valid),
    .io_enable_bits_taskID(const8_io_enable_bits_taskID),
    .io_Out_ready(const8_io_Out_ready),
    .io_Out_valid(const8_io_Out_valid),
    .io_Out_bits_taskID(const8_io_Out_bits_taskID)
  );
  ConstFastNode_9 const9 ( // @[extracted_function_conv.scala 446:22]
    .clock(const9_clock),
    .reset(const9_reset),
    .io_enable_ready(const9_io_enable_ready),
    .io_enable_valid(const9_io_enable_valid),
    .io_enable_bits_taskID(const9_io_enable_bits_taskID),
    .io_Out_ready(const9_io_Out_ready),
    .io_Out_valid(const9_io_Out_valid)
  );
  ConstFastNode_10 const10 ( // @[extracted_function_conv.scala 449:23]
    .clock(const10_clock),
    .reset(const10_reset),
    .io_enable_ready(const10_io_enable_ready),
    .io_enable_valid(const10_io_enable_valid),
    .io_enable_bits_taskID(const10_io_enable_bits_taskID),
    .io_Out_ready(const10_io_Out_ready),
    .io_Out_valid(const10_io_Out_valid)
  );
  ConstFastNode_11 const11 ( // @[extracted_function_conv.scala 452:23]
    .clock(const11_clock),
    .reset(const11_reset),
    .io_enable_ready(const11_io_enable_ready),
    .io_enable_valid(const11_io_enable_valid),
    .io_enable_bits_taskID(const11_io_enable_bits_taskID),
    .io_Out_ready(const11_io_Out_ready),
    .io_Out_valid(const11_io_Out_valid)
  );
  ConstFastNode_12 const12 ( // @[extracted_function_conv.scala 455:23]
    .clock(const12_clock),
    .reset(const12_reset),
    .io_enable_ready(const12_io_enable_ready),
    .io_enable_valid(const12_io_enable_valid),
    .io_enable_bits_taskID(const12_io_enable_bits_taskID),
    .io_Out_ready(const12_io_Out_ready),
    .io_Out_valid(const12_io_Out_valid)
  );
  ConstFastNode_13 const13 ( // @[extracted_function_conv.scala 458:23]
    .clock(const13_clock),
    .reset(const13_reset),
    .io_enable_ready(const13_io_enable_ready),
    .io_enable_valid(const13_io_enable_valid),
    .io_enable_bits_taskID(const13_io_enable_bits_taskID),
    .io_Out_ready(const13_io_Out_ready),
    .io_Out_valid(const13_io_Out_valid)
  );
  ConstFastNode_14 const14 ( // @[extracted_function_conv.scala 461:23]
    .clock(const14_clock),
    .reset(const14_reset),
    .io_enable_ready(const14_io_enable_ready),
    .io_enable_valid(const14_io_enable_valid),
    .io_enable_bits_taskID(const14_io_enable_bits_taskID),
    .io_Out_ready(const14_io_Out_ready),
    .io_Out_valid(const14_io_Out_valid)
  );
  ConstFastNode_15 const15 ( // @[extracted_function_conv.scala 464:23]
    .clock(const15_clock),
    .reset(const15_reset),
    .io_enable_ready(const15_io_enable_ready),
    .io_enable_valid(const15_io_enable_valid),
    .io_enable_bits_taskID(const15_io_enable_bits_taskID),
    .io_Out_ready(const15_io_Out_ready),
    .io_Out_valid(const15_io_Out_valid),
    .io_Out_bits_taskID(const15_io_Out_bits_taskID)
  );
  ConstFastNode_16 const16 ( // @[extracted_function_conv.scala 467:23]
    .clock(const16_clock),
    .reset(const16_reset),
    .io_enable_ready(const16_io_enable_ready),
    .io_enable_valid(const16_io_enable_valid),
    .io_enable_bits_taskID(const16_io_enable_bits_taskID),
    .io_Out_ready(const16_io_Out_ready),
    .io_Out_valid(const16_io_Out_valid)
  );
  ConstFastNode_17 const17 ( // @[extracted_function_conv.scala 470:23]
    .clock(const17_clock),
    .reset(const17_reset),
    .io_enable_ready(const17_io_enable_ready),
    .io_enable_valid(const17_io_enable_valid),
    .io_enable_bits_taskID(const17_io_enable_bits_taskID),
    .io_Out_ready(const17_io_Out_ready),
    .io_Out_valid(const17_io_Out_valid)
  );
  ConstFastNode_18 const18 ( // @[extracted_function_conv.scala 473:23]
    .clock(const18_clock),
    .reset(const18_reset),
    .io_enable_ready(const18_io_enable_ready),
    .io_enable_valid(const18_io_enable_valid),
    .io_enable_bits_taskID(const18_io_enable_bits_taskID),
    .io_Out_ready(const18_io_Out_ready),
    .io_Out_valid(const18_io_Out_valid)
  );
  ConstFastNode_19 const19 ( // @[extracted_function_conv.scala 476:23]
    .clock(const19_clock),
    .reset(const19_reset),
    .io_enable_ready(const19_io_enable_ready),
    .io_enable_valid(const19_io_enable_valid),
    .io_enable_bits_taskID(const19_io_enable_bits_taskID),
    .io_Out_ready(const19_io_Out_ready),
    .io_Out_valid(const19_io_Out_valid)
  );
  ConstFastNode_20 const20 ( // @[extracted_function_conv.scala 479:23]
    .clock(const20_clock),
    .reset(const20_reset),
    .io_enable_ready(const20_io_enable_ready),
    .io_enable_valid(const20_io_enable_valid),
    .io_enable_bits_taskID(const20_io_enable_bits_taskID),
    .io_Out_ready(const20_io_Out_ready),
    .io_Out_valid(const20_io_Out_valid)
  );
  ConstFastNode_21 const21 ( // @[extracted_function_conv.scala 482:23]
    .clock(const21_clock),
    .reset(const21_reset),
    .io_enable_ready(const21_io_enable_ready),
    .io_enable_valid(const21_io_enable_valid),
    .io_enable_bits_taskID(const21_io_enable_bits_taskID),
    .io_Out_ready(const21_io_Out_ready),
    .io_Out_valid(const21_io_Out_valid)
  );
  ConstFastNode_22 const22 ( // @[extracted_function_conv.scala 485:23]
    .clock(const22_clock),
    .reset(const22_reset),
    .io_enable_ready(const22_io_enable_ready),
    .io_enable_valid(const22_io_enable_valid),
    .io_enable_bits_taskID(const22_io_enable_bits_taskID),
    .io_Out_ready(const22_io_Out_ready),
    .io_Out_valid(const22_io_Out_valid)
  );
  ConstFastNode_23 const23 ( // @[extracted_function_conv.scala 488:23]
    .clock(const23_clock),
    .reset(const23_reset),
    .io_enable_ready(const23_io_enable_ready),
    .io_enable_valid(const23_io_enable_valid),
    .io_enable_bits_taskID(const23_io_enable_bits_taskID),
    .io_Out_ready(const23_io_Out_ready),
    .io_Out_valid(const23_io_Out_valid)
  );
  ConstFastNode_24 const24 ( // @[extracted_function_conv.scala 491:23]
    .clock(const24_clock),
    .reset(const24_reset),
    .io_enable_ready(const24_io_enable_ready),
    .io_enable_valid(const24_io_enable_valid),
    .io_enable_bits_taskID(const24_io_enable_bits_taskID),
    .io_Out_ready(const24_io_Out_ready),
    .io_Out_valid(const24_io_Out_valid)
  );
  ConstFastNode_25 const25 ( // @[extracted_function_conv.scala 494:23]
    .clock(const25_clock),
    .reset(const25_reset),
    .io_enable_ready(const25_io_enable_ready),
    .io_enable_valid(const25_io_enable_valid),
    .io_enable_bits_taskID(const25_io_enable_bits_taskID),
    .io_Out_ready(const25_io_Out_ready),
    .io_Out_valid(const25_io_Out_valid)
  );
  assign io_in_ready = InputSplitter_io_In_ready; // @[extracted_function_conv.scala 54:23]
  assign io_MemReq_valid = MemCtrl_io_MemReq_valid; // @[extracted_function_conv.scala 50:13]
  assign io_MemReq_bits_addr = MemCtrl_io_MemReq_bits_addr; // @[extracted_function_conv.scala 50:13]
  assign io_MemReq_bits_data = MemCtrl_io_MemReq_bits_data; // @[extracted_function_conv.scala 50:13]
  assign io_MemReq_bits_mask = MemCtrl_io_MemReq_bits_mask; // @[extracted_function_conv.scala 50:13]
  assign io_MemReq_bits_tag = MemCtrl_io_MemReq_bits_tag; // @[extracted_function_conv.scala 50:13]
  assign io_MemReq_bits_taskID = MemCtrl_io_MemReq_bits_taskID; // @[extracted_function_conv.scala 50:13]
  assign io_MemReq_bits_iswrite = MemCtrl_io_MemReq_bits_iswrite; // @[extracted_function_conv.scala 50:13]
  assign io_MemReq_bits_tile = 32'h0; // @[extracted_function_conv.scala 50:13]
  assign io_out_valid = ret_11_io_Out_valid; // @[extracted_function_conv.scala 1562:10]
  assign io_out_bits_enable_taskID = ret_11_io_Out_bits_enable_taskID; // @[extracted_function_conv.scala 1562:10]
  assign io_out_bits_enable_control = ret_11_io_Out_bits_enable_control; // @[extracted_function_conv.scala 1562:10]
  assign MemCtrl_clock = clock;
  assign MemCtrl_reset = reset;
  assign MemCtrl_io_WriteIn_0_valid = st_39_io_memReq_valid; // @[extracted_function_conv.scala 1128:25]
  assign MemCtrl_io_WriteIn_0_bits_address = st_39_io_memReq_bits_address; // @[extracted_function_conv.scala 1128:25]
  assign MemCtrl_io_WriteIn_0_bits_data = st_39_io_memReq_bits_data; // @[extracted_function_conv.scala 1128:25]
  assign MemCtrl_io_WriteIn_0_bits_taskID = st_39_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1128:25]
  assign MemCtrl_io_WriteIn_1_valid = st_47_io_memReq_valid; // @[extracted_function_conv.scala 1140:25]
  assign MemCtrl_io_WriteIn_1_bits_address = st_47_io_memReq_bits_address; // @[extracted_function_conv.scala 1140:25]
  assign MemCtrl_io_WriteIn_1_bits_data = st_47_io_memReq_bits_data; // @[extracted_function_conv.scala 1140:25]
  assign MemCtrl_io_WriteIn_1_bits_taskID = st_47_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1140:25]
  assign MemCtrl_io_WriteIn_2_valid = st_55_io_memReq_valid; // @[extracted_function_conv.scala 1152:25]
  assign MemCtrl_io_WriteIn_2_bits_address = st_55_io_memReq_bits_address; // @[extracted_function_conv.scala 1152:25]
  assign MemCtrl_io_WriteIn_2_bits_data = st_55_io_memReq_bits_data; // @[extracted_function_conv.scala 1152:25]
  assign MemCtrl_io_WriteIn_2_bits_taskID = st_55_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1152:25]
  assign MemCtrl_io_WriteIn_3_valid = st_64_io_memReq_valid; // @[extracted_function_conv.scala 1164:25]
  assign MemCtrl_io_WriteIn_3_bits_address = st_64_io_memReq_bits_address; // @[extracted_function_conv.scala 1164:25]
  assign MemCtrl_io_WriteIn_3_bits_data = st_64_io_memReq_bits_data; // @[extracted_function_conv.scala 1164:25]
  assign MemCtrl_io_WriteIn_3_bits_taskID = st_64_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1164:25]
  assign MemCtrl_io_WriteIn_4_valid = st_72_io_memReq_valid; // @[extracted_function_conv.scala 1176:25]
  assign MemCtrl_io_WriteIn_4_bits_address = st_72_io_memReq_bits_address; // @[extracted_function_conv.scala 1176:25]
  assign MemCtrl_io_WriteIn_4_bits_data = st_72_io_memReq_bits_data; // @[extracted_function_conv.scala 1176:25]
  assign MemCtrl_io_WriteIn_4_bits_taskID = st_72_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1176:25]
  assign MemCtrl_io_WriteIn_5_valid = st_80_io_memReq_valid; // @[extracted_function_conv.scala 1188:25]
  assign MemCtrl_io_WriteIn_5_bits_address = st_80_io_memReq_bits_address; // @[extracted_function_conv.scala 1188:25]
  assign MemCtrl_io_WriteIn_5_bits_data = st_80_io_memReq_bits_data; // @[extracted_function_conv.scala 1188:25]
  assign MemCtrl_io_WriteIn_5_bits_taskID = st_80_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1188:25]
  assign MemCtrl_io_WriteIn_6_valid = st_88_io_memReq_valid; // @[extracted_function_conv.scala 1200:25]
  assign MemCtrl_io_WriteIn_6_bits_address = st_88_io_memReq_bits_address; // @[extracted_function_conv.scala 1200:25]
  assign MemCtrl_io_WriteIn_6_bits_data = st_88_io_memReq_bits_data; // @[extracted_function_conv.scala 1200:25]
  assign MemCtrl_io_WriteIn_6_bits_taskID = st_88_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1200:25]
  assign MemCtrl_io_WriteIn_7_valid = st_96_io_memReq_valid; // @[extracted_function_conv.scala 1212:25]
  assign MemCtrl_io_WriteIn_7_bits_address = st_96_io_memReq_bits_address; // @[extracted_function_conv.scala 1212:25]
  assign MemCtrl_io_WriteIn_7_bits_data = st_96_io_memReq_bits_data; // @[extracted_function_conv.scala 1212:25]
  assign MemCtrl_io_WriteIn_7_bits_taskID = st_96_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1212:25]
  assign MemCtrl_io_WriteIn_8_valid = st_104_io_memReq_valid; // @[extracted_function_conv.scala 1224:25]
  assign MemCtrl_io_WriteIn_8_bits_address = st_104_io_memReq_bits_address; // @[extracted_function_conv.scala 1224:25]
  assign MemCtrl_io_WriteIn_8_bits_data = st_104_io_memReq_bits_data; // @[extracted_function_conv.scala 1224:25]
  assign MemCtrl_io_WriteIn_8_bits_taskID = st_104_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1224:25]
  assign MemCtrl_io_ReadIn_0_valid = ld_29_io_memReq_valid; // @[extracted_function_conv.scala 1116:24]
  assign MemCtrl_io_ReadIn_0_bits_address = ld_29_io_memReq_bits_address; // @[extracted_function_conv.scala 1116:24]
  assign MemCtrl_io_ReadIn_0_bits_taskID = ld_29_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1116:24]
  assign MemCtrl_io_ReadIn_1_valid = ld_30_io_memReq_valid; // @[extracted_function_conv.scala 1120:24]
  assign MemCtrl_io_ReadIn_1_bits_address = ld_30_io_memReq_bits_address; // @[extracted_function_conv.scala 1120:24]
  assign MemCtrl_io_ReadIn_1_bits_taskID = ld_30_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1120:24]
  assign MemCtrl_io_ReadIn_2_valid = ld_35_io_memReq_valid; // @[extracted_function_conv.scala 1124:24]
  assign MemCtrl_io_ReadIn_2_bits_address = ld_35_io_memReq_bits_address; // @[extracted_function_conv.scala 1124:24]
  assign MemCtrl_io_ReadIn_2_bits_taskID = ld_35_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1124:24]
  assign MemCtrl_io_ReadIn_3_valid = ld_40_io_memReq_valid; // @[extracted_function_conv.scala 1132:24]
  assign MemCtrl_io_ReadIn_3_bits_address = ld_40_io_memReq_bits_address; // @[extracted_function_conv.scala 1132:24]
  assign MemCtrl_io_ReadIn_3_bits_taskID = ld_40_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1132:24]
  assign MemCtrl_io_ReadIn_4_valid = ld_43_io_memReq_valid; // @[extracted_function_conv.scala 1136:24]
  assign MemCtrl_io_ReadIn_4_bits_address = ld_43_io_memReq_bits_address; // @[extracted_function_conv.scala 1136:24]
  assign MemCtrl_io_ReadIn_4_bits_taskID = ld_43_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1136:24]
  assign MemCtrl_io_ReadIn_5_valid = ld_48_io_memReq_valid; // @[extracted_function_conv.scala 1144:24]
  assign MemCtrl_io_ReadIn_5_bits_address = ld_48_io_memReq_bits_address; // @[extracted_function_conv.scala 1144:24]
  assign MemCtrl_io_ReadIn_5_bits_taskID = ld_48_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1144:24]
  assign MemCtrl_io_ReadIn_6_valid = ld_51_io_memReq_valid; // @[extracted_function_conv.scala 1148:24]
  assign MemCtrl_io_ReadIn_6_bits_address = ld_51_io_memReq_bits_address; // @[extracted_function_conv.scala 1148:24]
  assign MemCtrl_io_ReadIn_6_bits_taskID = ld_51_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1148:24]
  assign MemCtrl_io_ReadIn_7_valid = ld_56_io_memReq_valid; // @[extracted_function_conv.scala 1156:24]
  assign MemCtrl_io_ReadIn_7_bits_address = ld_56_io_memReq_bits_address; // @[extracted_function_conv.scala 1156:24]
  assign MemCtrl_io_ReadIn_7_bits_taskID = ld_56_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1156:24]
  assign MemCtrl_io_ReadIn_8_valid = ld_60_io_memReq_valid; // @[extracted_function_conv.scala 1160:24]
  assign MemCtrl_io_ReadIn_8_bits_address = ld_60_io_memReq_bits_address; // @[extracted_function_conv.scala 1160:24]
  assign MemCtrl_io_ReadIn_8_bits_taskID = ld_60_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1160:24]
  assign MemCtrl_io_ReadIn_9_valid = ld_65_io_memReq_valid; // @[extracted_function_conv.scala 1168:24]
  assign MemCtrl_io_ReadIn_9_bits_address = ld_65_io_memReq_bits_address; // @[extracted_function_conv.scala 1168:24]
  assign MemCtrl_io_ReadIn_9_bits_taskID = ld_65_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1168:24]
  assign MemCtrl_io_ReadIn_10_valid = ld_68_io_memReq_valid; // @[extracted_function_conv.scala 1172:25]
  assign MemCtrl_io_ReadIn_10_bits_address = ld_68_io_memReq_bits_address; // @[extracted_function_conv.scala 1172:25]
  assign MemCtrl_io_ReadIn_10_bits_taskID = ld_68_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1172:25]
  assign MemCtrl_io_ReadIn_11_valid = ld_73_io_memReq_valid; // @[extracted_function_conv.scala 1180:25]
  assign MemCtrl_io_ReadIn_11_bits_address = ld_73_io_memReq_bits_address; // @[extracted_function_conv.scala 1180:25]
  assign MemCtrl_io_ReadIn_11_bits_taskID = ld_73_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1180:25]
  assign MemCtrl_io_ReadIn_12_valid = ld_76_io_memReq_valid; // @[extracted_function_conv.scala 1184:25]
  assign MemCtrl_io_ReadIn_12_bits_address = ld_76_io_memReq_bits_address; // @[extracted_function_conv.scala 1184:25]
  assign MemCtrl_io_ReadIn_12_bits_taskID = ld_76_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1184:25]
  assign MemCtrl_io_ReadIn_13_valid = ld_81_io_memReq_valid; // @[extracted_function_conv.scala 1192:25]
  assign MemCtrl_io_ReadIn_13_bits_address = ld_81_io_memReq_bits_address; // @[extracted_function_conv.scala 1192:25]
  assign MemCtrl_io_ReadIn_13_bits_taskID = ld_81_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1192:25]
  assign MemCtrl_io_ReadIn_14_valid = ld_84_io_memReq_valid; // @[extracted_function_conv.scala 1196:25]
  assign MemCtrl_io_ReadIn_14_bits_address = ld_84_io_memReq_bits_address; // @[extracted_function_conv.scala 1196:25]
  assign MemCtrl_io_ReadIn_14_bits_taskID = ld_84_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1196:25]
  assign MemCtrl_io_ReadIn_15_valid = ld_89_io_memReq_valid; // @[extracted_function_conv.scala 1204:25]
  assign MemCtrl_io_ReadIn_15_bits_address = ld_89_io_memReq_bits_address; // @[extracted_function_conv.scala 1204:25]
  assign MemCtrl_io_ReadIn_15_bits_taskID = ld_89_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1204:25]
  assign MemCtrl_io_ReadIn_16_valid = ld_92_io_memReq_valid; // @[extracted_function_conv.scala 1208:25]
  assign MemCtrl_io_ReadIn_16_bits_address = ld_92_io_memReq_bits_address; // @[extracted_function_conv.scala 1208:25]
  assign MemCtrl_io_ReadIn_16_bits_taskID = ld_92_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1208:25]
  assign MemCtrl_io_ReadIn_17_valid = ld_97_io_memReq_valid; // @[extracted_function_conv.scala 1216:25]
  assign MemCtrl_io_ReadIn_17_bits_address = ld_97_io_memReq_bits_address; // @[extracted_function_conv.scala 1216:25]
  assign MemCtrl_io_ReadIn_17_bits_taskID = ld_97_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1216:25]
  assign MemCtrl_io_ReadIn_18_valid = ld_100_io_memReq_valid; // @[extracted_function_conv.scala 1220:25]
  assign MemCtrl_io_ReadIn_18_bits_address = ld_100_io_memReq_bits_address; // @[extracted_function_conv.scala 1220:25]
  assign MemCtrl_io_ReadIn_18_bits_taskID = ld_100_io_memReq_bits_taskID; // @[extracted_function_conv.scala 1220:25]
  assign MemCtrl_io_MemResp_valid = io_MemResp_valid; // @[extracted_function_conv.scala 51:22]
  assign MemCtrl_io_MemResp_bits_data = io_MemResp_bits_data; // @[extracted_function_conv.scala 51:22]
  assign MemCtrl_io_MemResp_bits_tag = io_MemResp_bits_tag; // @[extracted_function_conv.scala 51:22]
  assign MemCtrl_io_MemResp_bits_iswrite = io_MemResp_bits_iswrite; // @[extracted_function_conv.scala 51:22]
  assign MemCtrl_io_MemReq_ready = io_MemReq_ready; // @[extracted_function_conv.scala 50:13]
  assign InputSplitter_clock = clock;
  assign InputSplitter_reset = reset;
  assign InputSplitter_io_In_valid = io_in_valid; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_enable_taskID = io_in_bits_enable_taskID; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_enable_control = io_in_bits_enable_control; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field5_data = io_in_bits_data_field5_data; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field4_data = io_in_bits_data_field4_data; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field3_data = io_in_bits_data_field3_data; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field2_taskID = io_in_bits_data_field2_taskID; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field2_data = io_in_bits_data_field2_data; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field1_predicate = io_in_bits_data_field1_predicate; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field1_taskID = io_in_bits_data_field1_taskID; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field1_data = io_in_bits_data_field1_data; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field0_taskID = io_in_bits_data_field0_taskID; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_In_bits_data_field0_data = io_in_bits_data_field0_data; // @[extracted_function_conv.scala 54:23]
  assign InputSplitter_io_Out_enable_ready = bb_entry0_io_predicateIn_0_ready; // @[extracted_function_conv.scala 502:31]
  assign InputSplitter_io_Out_data_field5_0_ready = Loop_1_io_InLiveIn_0_ready; // @[extracted_function_conv.scala 590:25]
  assign InputSplitter_io_Out_data_field5_1_ready = binaryOp_mul0_io_LeftIO_ready; // @[extracted_function_conv.scala 1536:27]
  assign InputSplitter_io_Out_data_field4_0_ready = binaryOp_mul0_io_RightIO_ready; // @[extracted_function_conv.scala 1534:28]
  assign InputSplitter_io_Out_data_field3_0_ready = binaryOp_add1_io_RightIO_ready; // @[extracted_function_conv.scala 1532:28]
  assign InputSplitter_io_Out_data_field2_0_ready = Loop_1_io_InLiveIn_4_ready; // @[extracted_function_conv.scala 598:25]
  assign InputSplitter_io_Out_data_field1_0_ready = Loop_1_io_InLiveIn_3_ready; // @[extracted_function_conv.scala 596:25]
  assign InputSplitter_io_Out_data_field1_1_ready = Gep_arrayidx252_io_baseAddress_ready; // @[extracted_function_conv.scala 1516:34]
  assign InputSplitter_io_Out_data_field1_2_ready = Gep_arrayidx383_io_baseAddress_ready; // @[extracted_function_conv.scala 1518:34]
  assign InputSplitter_io_Out_data_field1_3_ready = Gep_arrayidx514_io_baseAddress_ready; // @[extracted_function_conv.scala 1520:34]
  assign InputSplitter_io_Out_data_field1_4_ready = Gep_arrayidx625_io_baseAddress_ready; // @[extracted_function_conv.scala 1522:34]
  assign InputSplitter_io_Out_data_field1_5_ready = Gep_arrayidx746_io_baseAddress_ready; // @[extracted_function_conv.scala 1524:34]
  assign InputSplitter_io_Out_data_field1_6_ready = Gep_arrayidx867_io_baseAddress_ready; // @[extracted_function_conv.scala 1526:34]
  assign InputSplitter_io_Out_data_field1_7_ready = Gep_arrayidx978_io_baseAddress_ready; // @[extracted_function_conv.scala 1528:34]
  assign InputSplitter_io_Out_data_field1_8_ready = Gep_arrayidx1099_io_baseAddress_ready; // @[extracted_function_conv.scala 1530:35]
  assign InputSplitter_io_Out_data_field0_0_ready = Loop_1_io_InLiveIn_2_ready; // @[extracted_function_conv.scala 594:25]
  assign Loop_0_clock = clock;
  assign Loop_0_reset = reset;
  assign Loop_0_io_enable_valid = br_22_io_Out_0_valid; // @[extracted_function_conv.scala 534:20]
  assign Loop_0_io_enable_bits_taskID = br_22_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 534:20]
  assign Loop_0_io_enable_bits_control = br_22_io_Out_0_bits_control; // @[extracted_function_conv.scala 534:20]
  assign Loop_0_io_InLiveIn_0_valid = binaryOp_mul821_io_Out_0_valid; // @[extracted_function_conv.scala 558:25]
  assign Loop_0_io_InLiveIn_0_bits_data = binaryOp_mul821_io_Out_0_bits_data; // @[extracted_function_conv.scala 558:25]
  assign Loop_0_io_InLiveIn_1_valid = binaryOp_mul720_io_Out_0_valid; // @[extracted_function_conv.scala 560:25]
  assign Loop_0_io_InLiveIn_1_bits_data = binaryOp_mul720_io_Out_0_bits_data; // @[extracted_function_conv.scala 560:25]
  assign Loop_0_io_InLiveIn_2_valid = binaryOp_sub16_io_Out_0_valid; // @[extracted_function_conv.scala 562:25]
  assign Loop_0_io_InLiveIn_2_bits_data = binaryOp_sub16_io_Out_0_bits_data; // @[extracted_function_conv.scala 562:25]
  assign Loop_0_io_InLiveIn_3_valid = binaryOp_sub619_io_Out_0_valid; // @[extracted_function_conv.scala 564:25]
  assign Loop_0_io_InLiveIn_3_bits_data = binaryOp_sub619_io_Out_0_bits_data; // @[extracted_function_conv.scala 564:25]
  assign Loop_0_io_InLiveIn_4_valid = Loop_1_io_OutLiveIn_field12_0_valid; // @[extracted_function_conv.scala 566:25]
  assign Loop_0_io_InLiveIn_4_bits_predicate = Loop_1_io_OutLiveIn_field12_0_bits_predicate; // @[extracted_function_conv.scala 566:25]
  assign Loop_0_io_InLiveIn_4_bits_taskID = Loop_1_io_OutLiveIn_field12_0_bits_taskID; // @[extracted_function_conv.scala 566:25]
  assign Loop_0_io_InLiveIn_4_bits_data = Loop_1_io_OutLiveIn_field12_0_bits_data; // @[extracted_function_conv.scala 566:25]
  assign Loop_0_io_InLiveIn_5_valid = Loop_1_io_OutLiveIn_field1_0_valid; // @[extracted_function_conv.scala 568:25]
  assign Loop_0_io_InLiveIn_5_bits_data = Loop_1_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_conv.scala 568:25]
  assign Loop_0_io_InLiveIn_6_valid = Loop_1_io_OutLiveIn_field9_0_valid; // @[extracted_function_conv.scala 570:25]
  assign Loop_0_io_InLiveIn_6_bits_predicate = Loop_1_io_OutLiveIn_field9_0_bits_predicate; // @[extracted_function_conv.scala 570:25]
  assign Loop_0_io_InLiveIn_6_bits_taskID = Loop_1_io_OutLiveIn_field9_0_bits_taskID; // @[extracted_function_conv.scala 570:25]
  assign Loop_0_io_InLiveIn_6_bits_data = Loop_1_io_OutLiveIn_field9_0_bits_data; // @[extracted_function_conv.scala 570:25]
  assign Loop_0_io_InLiveIn_7_valid = Loop_1_io_OutLiveIn_field8_0_valid; // @[extracted_function_conv.scala 572:25]
  assign Loop_0_io_InLiveIn_7_bits_predicate = Loop_1_io_OutLiveIn_field8_0_bits_predicate; // @[extracted_function_conv.scala 572:25]
  assign Loop_0_io_InLiveIn_7_bits_taskID = Loop_1_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_conv.scala 572:25]
  assign Loop_0_io_InLiveIn_7_bits_data = Loop_1_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_conv.scala 572:25]
  assign Loop_0_io_InLiveIn_8_valid = Loop_1_io_OutLiveIn_field7_0_valid; // @[extracted_function_conv.scala 574:25]
  assign Loop_0_io_InLiveIn_8_bits_predicate = Loop_1_io_OutLiveIn_field7_0_bits_predicate; // @[extracted_function_conv.scala 574:25]
  assign Loop_0_io_InLiveIn_8_bits_taskID = Loop_1_io_OutLiveIn_field7_0_bits_taskID; // @[extracted_function_conv.scala 574:25]
  assign Loop_0_io_InLiveIn_8_bits_data = Loop_1_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_conv.scala 574:25]
  assign Loop_0_io_InLiveIn_9_valid = Loop_1_io_OutLiveIn_field11_0_valid; // @[extracted_function_conv.scala 576:25]
  assign Loop_0_io_InLiveIn_9_bits_predicate = Loop_1_io_OutLiveIn_field11_0_bits_predicate; // @[extracted_function_conv.scala 576:25]
  assign Loop_0_io_InLiveIn_9_bits_taskID = Loop_1_io_OutLiveIn_field11_0_bits_taskID; // @[extracted_function_conv.scala 576:25]
  assign Loop_0_io_InLiveIn_9_bits_data = Loop_1_io_OutLiveIn_field11_0_bits_data; // @[extracted_function_conv.scala 576:25]
  assign Loop_0_io_InLiveIn_10_valid = Loop_1_io_OutLiveIn_field4_0_valid; // @[extracted_function_conv.scala 578:26]
  assign Loop_0_io_InLiveIn_10_bits_taskID = Loop_1_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_conv.scala 578:26]
  assign Loop_0_io_InLiveIn_10_bits_data = Loop_1_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_conv.scala 578:26]
  assign Loop_0_io_InLiveIn_11_valid = Loop_1_io_OutLiveIn_field2_0_valid; // @[extracted_function_conv.scala 580:26]
  assign Loop_0_io_InLiveIn_11_bits_taskID = Loop_1_io_OutLiveIn_field2_0_bits_taskID; // @[extracted_function_conv.scala 580:26]
  assign Loop_0_io_InLiveIn_11_bits_data = Loop_1_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_conv.scala 580:26]
  assign Loop_0_io_InLiveIn_12_valid = Loop_1_io_OutLiveIn_field6_0_valid; // @[extracted_function_conv.scala 582:26]
  assign Loop_0_io_InLiveIn_12_bits_predicate = Loop_1_io_OutLiveIn_field6_0_bits_predicate; // @[extracted_function_conv.scala 582:26]
  assign Loop_0_io_InLiveIn_12_bits_taskID = Loop_1_io_OutLiveIn_field6_0_bits_taskID; // @[extracted_function_conv.scala 582:26]
  assign Loop_0_io_InLiveIn_12_bits_data = Loop_1_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_conv.scala 582:26]
  assign Loop_0_io_InLiveIn_13_valid = Loop_1_io_OutLiveIn_field10_0_valid; // @[extracted_function_conv.scala 584:26]
  assign Loop_0_io_InLiveIn_13_bits_predicate = Loop_1_io_OutLiveIn_field10_0_bits_predicate; // @[extracted_function_conv.scala 584:26]
  assign Loop_0_io_InLiveIn_13_bits_taskID = Loop_1_io_OutLiveIn_field10_0_bits_taskID; // @[extracted_function_conv.scala 584:26]
  assign Loop_0_io_InLiveIn_13_bits_data = Loop_1_io_OutLiveIn_field10_0_bits_data; // @[extracted_function_conv.scala 584:26]
  assign Loop_0_io_InLiveIn_14_valid = Loop_1_io_OutLiveIn_field3_0_valid; // @[extracted_function_conv.scala 586:26]
  assign Loop_0_io_InLiveIn_14_bits_predicate = Loop_1_io_OutLiveIn_field3_0_bits_predicate; // @[extracted_function_conv.scala 586:26]
  assign Loop_0_io_InLiveIn_14_bits_taskID = Loop_1_io_OutLiveIn_field3_0_bits_taskID; // @[extracted_function_conv.scala 586:26]
  assign Loop_0_io_InLiveIn_14_bits_data = Loop_1_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_conv.scala 586:26]
  assign Loop_0_io_InLiveIn_15_valid = Loop_1_io_OutLiveIn_field5_0_valid; // @[extracted_function_conv.scala 588:26]
  assign Loop_0_io_InLiveIn_15_bits_predicate = Loop_1_io_OutLiveIn_field5_0_bits_predicate; // @[extracted_function_conv.scala 588:26]
  assign Loop_0_io_InLiveIn_15_bits_taskID = Loop_1_io_OutLiveIn_field5_0_bits_taskID; // @[extracted_function_conv.scala 588:26]
  assign Loop_0_io_InLiveIn_15_bits_data = Loop_1_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_conv.scala 588:26]
  assign Loop_0_io_OutLiveIn_field15_0_ready = ld_40_io_GepAddr_ready; // @[extracted_function_conv.scala 668:20]
  assign Loop_0_io_OutLiveIn_field14_0_ready = ld_30_io_GepAddr_ready; // @[extracted_function_conv.scala 666:20]
  assign Loop_0_io_OutLiveIn_field13_0_ready = ld_81_io_GepAddr_ready; // @[extracted_function_conv.scala 664:20]
  assign Loop_0_io_OutLiveIn_field12_0_ready = ld_48_io_GepAddr_ready; // @[extracted_function_conv.scala 662:20]
  assign Loop_0_io_OutLiveIn_field11_0_ready = Gep_arrayidx28_io_baseAddress_ready; // @[extracted_function_conv.scala 660:33]
  assign Loop_0_io_OutLiveIn_field10_0_ready = Gep_arrayidx1834_io_baseAddress_ready; // @[extracted_function_conv.scala 642:35]
  assign Loop_0_io_OutLiveIn_field10_1_ready = Gep_arrayidx3042_io_baseAddress_ready; // @[extracted_function_conv.scala 644:35]
  assign Loop_0_io_OutLiveIn_field10_2_ready = Gep_arrayidx4350_io_baseAddress_ready; // @[extracted_function_conv.scala 646:35]
  assign Loop_0_io_OutLiveIn_field10_3_ready = Gep_arrayidx5459_io_baseAddress_ready; // @[extracted_function_conv.scala 648:35]
  assign Loop_0_io_OutLiveIn_field10_4_ready = Gep_arrayidx6667_io_baseAddress_ready; // @[extracted_function_conv.scala 650:35]
  assign Loop_0_io_OutLiveIn_field10_5_ready = Gep_arrayidx7875_io_baseAddress_ready; // @[extracted_function_conv.scala 652:35]
  assign Loop_0_io_OutLiveIn_field10_6_ready = Gep_arrayidx8983_io_baseAddress_ready; // @[extracted_function_conv.scala 654:35]
  assign Loop_0_io_OutLiveIn_field10_7_ready = Gep_arrayidx10191_io_baseAddress_ready; // @[extracted_function_conv.scala 656:36]
  assign Loop_0_io_OutLiveIn_field10_8_ready = Gep_arrayidx11399_io_baseAddress_ready; // @[extracted_function_conv.scala 658:36]
  assign Loop_0_io_OutLiveIn_field9_0_ready = ld_89_io_GepAddr_ready; // @[extracted_function_conv.scala 640:20]
  assign Loop_0_io_OutLiveIn_field8_0_ready = ld_56_io_GepAddr_ready; // @[extracted_function_conv.scala 638:20]
  assign Loop_0_io_OutLiveIn_field7_0_ready = ld_65_io_GepAddr_ready; // @[extracted_function_conv.scala 636:20]
  assign Loop_0_io_OutLiveIn_field6_0_ready = ld_73_io_GepAddr_ready; // @[extracted_function_conv.scala 634:20]
  assign Loop_0_io_OutLiveIn_field5_0_ready = binaryOp_sub1733_io_RightIO_ready; // @[extracted_function_conv.scala 632:31]
  assign Loop_0_io_OutLiveIn_field4_0_ready = ld_97_io_GepAddr_ready; // @[extracted_function_conv.scala 630:20]
  assign Loop_0_io_OutLiveIn_field3_0_ready = binaryOp_add8882_io_RightIO_ready; // @[extracted_function_conv.scala 628:31]
  assign Loop_0_io_OutLiveIn_field2_0_ready = binaryOp_add5358_io_RightIO_ready; // @[extracted_function_conv.scala 626:31]
  assign Loop_0_io_OutLiveIn_field1_0_ready = binaryOp_add1531_io_RightIO_ready; // @[extracted_function_conv.scala 624:31]
  assign Loop_0_io_OutLiveIn_field0_0_ready = binaryOp_add1327_io_RightIO_ready; // @[extracted_function_conv.scala 622:31]
  assign Loop_0_io_activate_loop_start_ready = bb_for_body124_io_predicateIn_1_ready; // @[extracted_function_conv.scala 518:36]
  assign Loop_0_io_activate_loop_back_ready = bb_for_body124_io_predicateIn_0_ready; // @[extracted_function_conv.scala 520:36]
  assign Loop_0_io_loopBack_0_valid = br_107_io_FalseOutput_0_valid; // @[extracted_function_conv.scala 536:25]
  assign Loop_0_io_loopBack_0_bits_taskID = br_107_io_FalseOutput_0_bits_taskID; // @[extracted_function_conv.scala 536:25]
  assign Loop_0_io_loopBack_0_bits_control = br_107_io_FalseOutput_0_bits_control; // @[extracted_function_conv.scala 536:25]
  assign Loop_0_io_loopFinish_0_valid = br_107_io_TrueOutput_0_valid; // @[extracted_function_conv.scala 538:27]
  assign Loop_0_io_loopFinish_0_bits_control = br_107_io_TrueOutput_0_bits_control; // @[extracted_function_conv.scala 538:27]
  assign Loop_0_io_CarryDepenIn_0_valid = binaryOp_inc105_io_Out_0_valid; // @[extracted_function_conv.scala 698:29]
  assign Loop_0_io_CarryDepenIn_0_bits_taskID = binaryOp_inc105_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 698:29]
  assign Loop_0_io_CarryDepenIn_0_bits_data = binaryOp_inc105_io_Out_0_bits_data; // @[extracted_function_conv.scala 698:29]
  assign Loop_0_io_CarryDepenOut_field0_0_ready = phi_conv_s1_x_031226_io_InData_1_ready; // @[extracted_function_conv.scala 708:37]
  assign Loop_0_io_loopExit_0_ready = bb_for_cond_cleanup113_io_predicateIn_0_ready; // @[extracted_function_conv.scala 516:44]
  assign Loop_1_clock = clock;
  assign Loop_1_reset = reset;
  assign Loop_1_io_enable_valid = br_10_io_Out_0_valid; // @[extracted_function_conv.scala 540:20]
  assign Loop_1_io_enable_bits_taskID = br_10_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 540:20]
  assign Loop_1_io_enable_bits_control = br_10_io_Out_0_bits_control; // @[extracted_function_conv.scala 540:20]
  assign Loop_1_io_InLiveIn_0_valid = InputSplitter_io_Out_data_field5_0_valid; // @[extracted_function_conv.scala 590:25]
  assign Loop_1_io_InLiveIn_0_bits_data = InputSplitter_io_Out_data_field5_0_bits_data; // @[extracted_function_conv.scala 590:25]
  assign Loop_1_io_InLiveIn_1_valid = binaryOp_add1_io_Out_0_valid; // @[extracted_function_conv.scala 592:25]
  assign Loop_1_io_InLiveIn_1_bits_data = binaryOp_add1_io_Out_0_bits_data; // @[extracted_function_conv.scala 592:25]
  assign Loop_1_io_InLiveIn_2_valid = InputSplitter_io_Out_data_field0_0_valid; // @[extracted_function_conv.scala 594:25]
  assign Loop_1_io_InLiveIn_2_bits_taskID = InputSplitter_io_Out_data_field0_0_bits_taskID; // @[extracted_function_conv.scala 594:25]
  assign Loop_1_io_InLiveIn_2_bits_data = InputSplitter_io_Out_data_field0_0_bits_data; // @[extracted_function_conv.scala 594:25]
  assign Loop_1_io_InLiveIn_3_valid = InputSplitter_io_Out_data_field1_0_valid; // @[extracted_function_conv.scala 596:25]
  assign Loop_1_io_InLiveIn_3_bits_predicate = InputSplitter_io_Out_data_field1_0_bits_predicate; // @[extracted_function_conv.scala 596:25]
  assign Loop_1_io_InLiveIn_3_bits_taskID = InputSplitter_io_Out_data_field1_0_bits_taskID; // @[extracted_function_conv.scala 596:25]
  assign Loop_1_io_InLiveIn_3_bits_data = InputSplitter_io_Out_data_field1_0_bits_data; // @[extracted_function_conv.scala 596:25]
  assign Loop_1_io_InLiveIn_4_valid = InputSplitter_io_Out_data_field2_0_valid; // @[extracted_function_conv.scala 598:25]
  assign Loop_1_io_InLiveIn_4_bits_taskID = InputSplitter_io_Out_data_field2_0_bits_taskID; // @[extracted_function_conv.scala 598:25]
  assign Loop_1_io_InLiveIn_4_bits_data = InputSplitter_io_Out_data_field2_0_bits_data; // @[extracted_function_conv.scala 598:25]
  assign Loop_1_io_InLiveIn_5_valid = Gep_arrayidx252_io_Out_0_valid; // @[extracted_function_conv.scala 600:25]
  assign Loop_1_io_InLiveIn_5_bits_predicate = Gep_arrayidx252_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 600:25]
  assign Loop_1_io_InLiveIn_5_bits_taskID = Gep_arrayidx252_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 600:25]
  assign Loop_1_io_InLiveIn_5_bits_data = Gep_arrayidx252_io_Out_0_bits_data; // @[extracted_function_conv.scala 600:25]
  assign Loop_1_io_InLiveIn_6_valid = Gep_arrayidx383_io_Out_0_valid; // @[extracted_function_conv.scala 602:25]
  assign Loop_1_io_InLiveIn_6_bits_predicate = Gep_arrayidx383_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 602:25]
  assign Loop_1_io_InLiveIn_6_bits_taskID = Gep_arrayidx383_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 602:25]
  assign Loop_1_io_InLiveIn_6_bits_data = Gep_arrayidx383_io_Out_0_bits_data; // @[extracted_function_conv.scala 602:25]
  assign Loop_1_io_InLiveIn_7_valid = Gep_arrayidx514_io_Out_0_valid; // @[extracted_function_conv.scala 604:25]
  assign Loop_1_io_InLiveIn_7_bits_predicate = Gep_arrayidx514_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 604:25]
  assign Loop_1_io_InLiveIn_7_bits_taskID = Gep_arrayidx514_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 604:25]
  assign Loop_1_io_InLiveIn_7_bits_data = Gep_arrayidx514_io_Out_0_bits_data; // @[extracted_function_conv.scala 604:25]
  assign Loop_1_io_InLiveIn_8_valid = Gep_arrayidx625_io_Out_0_valid; // @[extracted_function_conv.scala 606:25]
  assign Loop_1_io_InLiveIn_8_bits_predicate = Gep_arrayidx625_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 606:25]
  assign Loop_1_io_InLiveIn_8_bits_taskID = Gep_arrayidx625_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 606:25]
  assign Loop_1_io_InLiveIn_8_bits_data = Gep_arrayidx625_io_Out_0_bits_data; // @[extracted_function_conv.scala 606:25]
  assign Loop_1_io_InLiveIn_9_valid = Gep_arrayidx746_io_Out_0_valid; // @[extracted_function_conv.scala 608:25]
  assign Loop_1_io_InLiveIn_9_bits_predicate = Gep_arrayidx746_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 608:25]
  assign Loop_1_io_InLiveIn_9_bits_taskID = Gep_arrayidx746_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 608:25]
  assign Loop_1_io_InLiveIn_9_bits_data = Gep_arrayidx746_io_Out_0_bits_data; // @[extracted_function_conv.scala 608:25]
  assign Loop_1_io_InLiveIn_10_valid = Gep_arrayidx867_io_Out_0_valid; // @[extracted_function_conv.scala 610:26]
  assign Loop_1_io_InLiveIn_10_bits_predicate = Gep_arrayidx867_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 610:26]
  assign Loop_1_io_InLiveIn_10_bits_taskID = Gep_arrayidx867_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 610:26]
  assign Loop_1_io_InLiveIn_10_bits_data = Gep_arrayidx867_io_Out_0_bits_data; // @[extracted_function_conv.scala 610:26]
  assign Loop_1_io_InLiveIn_11_valid = Gep_arrayidx978_io_Out_0_valid; // @[extracted_function_conv.scala 612:26]
  assign Loop_1_io_InLiveIn_11_bits_predicate = Gep_arrayidx978_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 612:26]
  assign Loop_1_io_InLiveIn_11_bits_taskID = Gep_arrayidx978_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 612:26]
  assign Loop_1_io_InLiveIn_11_bits_data = Gep_arrayidx978_io_Out_0_bits_data; // @[extracted_function_conv.scala 612:26]
  assign Loop_1_io_InLiveIn_12_valid = Gep_arrayidx1099_io_Out_0_valid; // @[extracted_function_conv.scala 614:26]
  assign Loop_1_io_InLiveIn_12_bits_predicate = Gep_arrayidx1099_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 614:26]
  assign Loop_1_io_InLiveIn_12_bits_taskID = Gep_arrayidx1099_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 614:26]
  assign Loop_1_io_InLiveIn_12_bits_data = Gep_arrayidx1099_io_Out_0_bits_data; // @[extracted_function_conv.scala 614:26]
  assign Loop_1_io_OutLiveIn_field12_0_ready = Loop_0_io_InLiveIn_4_ready; // @[extracted_function_conv.scala 566:25]
  assign Loop_1_io_OutLiveIn_field11_0_ready = Loop_0_io_InLiveIn_9_ready; // @[extracted_function_conv.scala 576:25]
  assign Loop_1_io_OutLiveIn_field10_0_ready = Loop_0_io_InLiveIn_13_ready; // @[extracted_function_conv.scala 584:26]
  assign Loop_1_io_OutLiveIn_field9_0_ready = Loop_0_io_InLiveIn_6_ready; // @[extracted_function_conv.scala 570:25]
  assign Loop_1_io_OutLiveIn_field8_0_ready = Loop_0_io_InLiveIn_7_ready; // @[extracted_function_conv.scala 572:25]
  assign Loop_1_io_OutLiveIn_field7_0_ready = Loop_0_io_InLiveIn_8_ready; // @[extracted_function_conv.scala 574:25]
  assign Loop_1_io_OutLiveIn_field6_0_ready = Loop_0_io_InLiveIn_12_ready; // @[extracted_function_conv.scala 582:26]
  assign Loop_1_io_OutLiveIn_field5_0_ready = Loop_0_io_InLiveIn_15_ready; // @[extracted_function_conv.scala 588:26]
  assign Loop_1_io_OutLiveIn_field4_0_ready = Loop_0_io_InLiveIn_10_ready; // @[extracted_function_conv.scala 578:26]
  assign Loop_1_io_OutLiveIn_field3_0_ready = Loop_0_io_InLiveIn_14_ready; // @[extracted_function_conv.scala 586:26]
  assign Loop_1_io_OutLiveIn_field2_0_ready = Loop_0_io_InLiveIn_11_ready; // @[extracted_function_conv.scala 580:26]
  assign Loop_1_io_OutLiveIn_field1_0_ready = Loop_0_io_InLiveIn_5_ready; // @[extracted_function_conv.scala 568:25]
  assign Loop_1_io_OutLiveIn_field1_1_ready = binaryOp_sub16_io_RightIO_ready; // @[extracted_function_conv.scala 676:29]
  assign Loop_1_io_OutLiveIn_field1_2_ready = binaryOp_sub619_io_RightIO_ready; // @[extracted_function_conv.scala 678:30]
  assign Loop_1_io_OutLiveIn_field0_0_ready = binaryOp_mul315_io_RightIO_ready; // @[extracted_function_conv.scala 670:30]
  assign Loop_1_io_OutLiveIn_field0_1_ready = binaryOp_mul518_io_RightIO_ready; // @[extracted_function_conv.scala 672:30]
  assign Loop_1_io_OutLiveIn_field0_2_ready = binaryOp_mul720_io_RightIO_ready; // @[extracted_function_conv.scala 674:30]
  assign Loop_1_io_activate_loop_start_ready = bb_for_body2_io_predicateIn_1_ready; // @[extracted_function_conv.scala 512:34]
  assign Loop_1_io_activate_loop_back_ready = bb_for_body2_io_predicateIn_0_ready; // @[extracted_function_conv.scala 514:34]
  assign Loop_1_io_loopBack_0_valid = br_25_io_FalseOutput_0_valid; // @[extracted_function_conv.scala 542:25]
  assign Loop_1_io_loopBack_0_bits_taskID = br_25_io_FalseOutput_0_bits_taskID; // @[extracted_function_conv.scala 542:25]
  assign Loop_1_io_loopBack_0_bits_control = br_25_io_FalseOutput_0_bits_control; // @[extracted_function_conv.scala 542:25]
  assign Loop_1_io_loopFinish_0_valid = br_25_io_TrueOutput_0_valid; // @[extracted_function_conv.scala 544:27]
  assign Loop_1_io_loopFinish_0_bits_control = br_25_io_TrueOutput_0_bits_control; // @[extracted_function_conv.scala 544:27]
  assign Loop_1_io_CarryDepenIn_0_valid = binaryOp_inc12023_io_Out_0_valid; // @[extracted_function_conv.scala 700:29]
  assign Loop_1_io_CarryDepenIn_0_bits_taskID = binaryOp_inc12023_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 700:29]
  assign Loop_1_io_CarryDepenIn_0_bits_data = binaryOp_inc12023_io_Out_0_bits_data; // @[extracted_function_conv.scala 700:29]
  assign Loop_1_io_CarryDepenOut_field0_0_ready = phi_conv_s1_y_031312_io_InData_1_ready; // @[extracted_function_conv.scala 710:37]
  assign Loop_1_io_loopExit_0_ready = bb_for_cond_cleanup1_io_predicateIn_0_ready; // @[extracted_function_conv.scala 510:42]
  assign bb_entry0_clock = clock;
  assign bb_entry0_reset = reset;
  assign bb_entry0_io_predicateIn_0_valid = InputSplitter_io_Out_enable_valid; // @[extracted_function_conv.scala 502:31]
  assign bb_entry0_io_predicateIn_0_bits_taskID = InputSplitter_io_Out_enable_bits_taskID; // @[extracted_function_conv.scala 502:31]
  assign bb_entry0_io_predicateIn_0_bits_control = InputSplitter_io_Out_enable_bits_control; // @[extracted_function_conv.scala 502:31]
  assign bb_entry0_io_Out_0_ready = const0_io_enable_ready; // @[extracted_function_conv.scala 718:20]
  assign bb_entry0_io_Out_1_ready = const1_io_enable_ready; // @[extracted_function_conv.scala 720:20]
  assign bb_entry0_io_Out_2_ready = const2_io_enable_ready; // @[extracted_function_conv.scala 722:20]
  assign bb_entry0_io_Out_3_ready = const3_io_enable_ready; // @[extracted_function_conv.scala 724:20]
  assign bb_entry0_io_Out_4_ready = const4_io_enable_ready; // @[extracted_function_conv.scala 726:20]
  assign bb_entry0_io_Out_5_ready = const5_io_enable_ready; // @[extracted_function_conv.scala 728:20]
  assign bb_entry0_io_Out_6_ready = const6_io_enable_ready; // @[extracted_function_conv.scala 730:20]
  assign bb_entry0_io_Out_7_ready = const7_io_enable_ready; // @[extracted_function_conv.scala 732:20]
  assign bb_entry0_io_Out_8_ready = binaryOp_mul0_io_enable_ready; // @[extracted_function_conv.scala 734:27]
  assign bb_entry0_io_Out_9_ready = binaryOp_add1_io_enable_ready; // @[extracted_function_conv.scala 737:27]
  assign bb_entry0_io_Out_10_ready = Gep_arrayidx252_io_enable_ready; // @[extracted_function_conv.scala 740:29]
  assign bb_entry0_io_Out_11_ready = Gep_arrayidx383_io_enable_ready; // @[extracted_function_conv.scala 743:29]
  assign bb_entry0_io_Out_12_ready = Gep_arrayidx514_io_enable_ready; // @[extracted_function_conv.scala 746:29]
  assign bb_entry0_io_Out_13_ready = Gep_arrayidx625_io_enable_ready; // @[extracted_function_conv.scala 749:29]
  assign bb_entry0_io_Out_14_ready = Gep_arrayidx746_io_enable_ready; // @[extracted_function_conv.scala 752:29]
  assign bb_entry0_io_Out_15_ready = Gep_arrayidx867_io_enable_ready; // @[extracted_function_conv.scala 755:29]
  assign bb_entry0_io_Out_16_ready = Gep_arrayidx978_io_enable_ready; // @[extracted_function_conv.scala 758:29]
  assign bb_entry0_io_Out_17_ready = Gep_arrayidx1099_io_enable_ready; // @[extracted_function_conv.scala 761:30]
  assign bb_entry0_io_Out_18_ready = br_10_io_enable_ready; // @[extracted_function_conv.scala 764:19]
  assign bb_for_cond_cleanup1_clock = clock;
  assign bb_for_cond_cleanup1_reset = reset;
  assign bb_for_cond_cleanup1_io_predicateIn_0_valid = Loop_1_io_loopExit_0_valid; // @[extracted_function_conv.scala 510:42]
  assign bb_for_cond_cleanup1_io_predicateIn_0_bits_taskID = Loop_1_io_loopExit_0_bits_taskID; // @[extracted_function_conv.scala 510:42]
  assign bb_for_cond_cleanup1_io_predicateIn_0_bits_control = Loop_1_io_loopExit_0_bits_control; // @[extracted_function_conv.scala 510:42]
  assign bb_for_cond_cleanup1_io_Out_0_ready = ret_11_io_In_enable_ready; // @[extracted_function_conv.scala 767:23]
  assign bb_for_body2_clock = clock;
  assign bb_for_body2_reset = reset;
  assign bb_for_body2_io_MaskBB_0_ready = phi_conv_s1_y_031312_io_Mask_ready; // @[extracted_function_conv.scala 1100:32]
  assign bb_for_body2_io_Out_0_ready = const8_io_enable_ready; // @[extracted_function_conv.scala 770:20]
  assign bb_for_body2_io_Out_1_ready = const9_io_enable_ready; // @[extracted_function_conv.scala 772:20]
  assign bb_for_body2_io_Out_2_ready = const10_io_enable_ready; // @[extracted_function_conv.scala 774:21]
  assign bb_for_body2_io_Out_3_ready = const11_io_enable_ready; // @[extracted_function_conv.scala 776:21]
  assign bb_for_body2_io_Out_4_ready = const12_io_enable_ready; // @[extracted_function_conv.scala 778:21]
  assign bb_for_body2_io_Out_5_ready = phi_conv_s1_y_031312_io_enable_ready; // @[extracted_function_conv.scala 780:34]
  assign bb_for_body2_io_Out_6_ready = binaryOp_mul113_io_enable_ready; // @[extracted_function_conv.scala 783:29]
  assign bb_for_body2_io_Out_7_ready = binaryOp_add214_io_enable_ready; // @[extracted_function_conv.scala 786:29]
  assign bb_for_body2_io_Out_8_ready = binaryOp_mul315_io_enable_ready; // @[extracted_function_conv.scala 789:29]
  assign bb_for_body2_io_Out_9_ready = binaryOp_sub16_io_enable_ready; // @[extracted_function_conv.scala 792:28]
  assign bb_for_body2_io_Out_10_ready = binaryOp_add417_io_enable_ready; // @[extracted_function_conv.scala 795:29]
  assign bb_for_body2_io_Out_11_ready = binaryOp_mul518_io_enable_ready; // @[extracted_function_conv.scala 798:29]
  assign bb_for_body2_io_Out_12_ready = binaryOp_sub619_io_enable_ready; // @[extracted_function_conv.scala 801:29]
  assign bb_for_body2_io_Out_13_ready = binaryOp_mul720_io_enable_ready; // @[extracted_function_conv.scala 804:29]
  assign bb_for_body2_io_Out_14_ready = binaryOp_mul821_io_enable_ready; // @[extracted_function_conv.scala 807:29]
  assign bb_for_body2_io_Out_15_ready = br_22_io_enable_ready; // @[extracted_function_conv.scala 810:19]
  assign bb_for_body2_io_predicateIn_0_valid = Loop_1_io_activate_loop_back_valid; // @[extracted_function_conv.scala 514:34]
  assign bb_for_body2_io_predicateIn_0_bits_taskID = Loop_1_io_activate_loop_back_bits_taskID; // @[extracted_function_conv.scala 514:34]
  assign bb_for_body2_io_predicateIn_0_bits_control = Loop_1_io_activate_loop_back_bits_control; // @[extracted_function_conv.scala 514:34]
  assign bb_for_body2_io_predicateIn_1_valid = Loop_1_io_activate_loop_start_valid; // @[extracted_function_conv.scala 512:34]
  assign bb_for_body2_io_predicateIn_1_bits_taskID = Loop_1_io_activate_loop_start_bits_taskID; // @[extracted_function_conv.scala 512:34]
  assign bb_for_body2_io_predicateIn_1_bits_control = Loop_1_io_activate_loop_start_bits_control; // @[extracted_function_conv.scala 512:34]
  assign bb_for_cond_cleanup113_clock = clock;
  assign bb_for_cond_cleanup113_reset = reset;
  assign bb_for_cond_cleanup113_io_predicateIn_0_valid = Loop_0_io_loopExit_0_valid; // @[extracted_function_conv.scala 516:44]
  assign bb_for_cond_cleanup113_io_predicateIn_0_bits_taskID = Loop_0_io_loopExit_0_bits_taskID; // @[extracted_function_conv.scala 516:44]
  assign bb_for_cond_cleanup113_io_predicateIn_0_bits_control = Loop_0_io_loopExit_0_bits_control; // @[extracted_function_conv.scala 516:44]
  assign bb_for_cond_cleanup113_io_Out_0_ready = const13_io_enable_ready; // @[extracted_function_conv.scala 813:21]
  assign bb_for_cond_cleanup113_io_Out_1_ready = const14_io_enable_ready; // @[extracted_function_conv.scala 815:21]
  assign bb_for_cond_cleanup113_io_Out_2_ready = binaryOp_inc12023_io_enable_ready; // @[extracted_function_conv.scala 817:31]
  assign bb_for_cond_cleanup113_io_Out_3_ready = icmp_exitcond31424_io_enable_ready; // @[extracted_function_conv.scala 820:32]
  assign bb_for_cond_cleanup113_io_Out_4_ready = br_25_io_enable_ready; // @[extracted_function_conv.scala 823:19]
  assign bb_for_body124_clock = clock;
  assign bb_for_body124_reset = reset;
  assign bb_for_body124_io_MaskBB_0_ready = phi_conv_s1_x_031226_io_Mask_ready; // @[extracted_function_conv.scala 1102:32]
  assign bb_for_body124_io_Out_0_ready = const15_io_enable_ready; // @[extracted_function_conv.scala 826:21]
  assign bb_for_body124_io_Out_1_ready = const16_io_enable_ready; // @[extracted_function_conv.scala 828:21]
  assign bb_for_body124_io_Out_2_ready = const17_io_enable_ready; // @[extracted_function_conv.scala 830:21]
  assign bb_for_body124_io_Out_3_ready = const18_io_enable_ready; // @[extracted_function_conv.scala 832:21]
  assign bb_for_body124_io_Out_4_ready = const19_io_enable_ready; // @[extracted_function_conv.scala 834:21]
  assign bb_for_body124_io_Out_5_ready = const20_io_enable_ready; // @[extracted_function_conv.scala 836:21]
  assign bb_for_body124_io_Out_6_ready = const21_io_enable_ready; // @[extracted_function_conv.scala 838:21]
  assign bb_for_body124_io_Out_7_ready = const22_io_enable_ready; // @[extracted_function_conv.scala 840:21]
  assign bb_for_body124_io_Out_8_ready = const23_io_enable_ready; // @[extracted_function_conv.scala 842:21]
  assign bb_for_body124_io_Out_9_ready = const24_io_enable_ready; // @[extracted_function_conv.scala 844:21]
  assign bb_for_body124_io_Out_10_ready = const25_io_enable_ready; // @[extracted_function_conv.scala 846:21]
  assign bb_for_body124_io_Out_11_ready = phi_conv_s1_x_031226_io_enable_ready; // @[extracted_function_conv.scala 848:34]
  assign bb_for_body124_io_Out_12_ready = binaryOp_add1327_io_enable_ready; // @[extracted_function_conv.scala 851:30]
  assign bb_for_body124_io_Out_13_ready = Gep_arrayidx28_io_enable_ready; // @[extracted_function_conv.scala 854:28]
  assign bb_for_body124_io_Out_14_ready = ld_29_io_enable_ready; // @[extracted_function_conv.scala 857:19]
  assign bb_for_body124_io_Out_15_ready = ld_30_io_enable_ready; // @[extracted_function_conv.scala 860:19]
  assign bb_for_body124_io_Out_16_ready = binaryOp_add1531_io_enable_ready; // @[extracted_function_conv.scala 863:30]
  assign bb_for_body124_io_Out_17_ready = binaryOp_mul1632_io_enable_ready; // @[extracted_function_conv.scala 866:30]
  assign bb_for_body124_io_Out_18_ready = binaryOp_sub1733_io_enable_ready; // @[extracted_function_conv.scala 869:30]
  assign bb_for_body124_io_Out_19_ready = Gep_arrayidx1834_io_enable_ready; // @[extracted_function_conv.scala 872:30]
  assign bb_for_body124_io_Out_20_ready = ld_35_io_enable_ready; // @[extracted_function_conv.scala 875:19]
  assign bb_for_body124_io_Out_21_ready = sextconv1936_io_enable_ready; // @[extracted_function_conv.scala 878:26]
  assign bb_for_body124_io_Out_22_ready = binaryOp_mul2037_io_enable_ready; // @[extracted_function_conv.scala 881:30]
  assign bb_for_body124_io_Out_23_ready = binaryOp_add2138_io_enable_ready; // @[extracted_function_conv.scala 884:30]
  assign bb_for_body124_io_Out_24_ready = st_39_io_enable_ready; // @[extracted_function_conv.scala 887:19]
  assign bb_for_body124_io_Out_25_ready = ld_40_io_enable_ready; // @[extracted_function_conv.scala 890:19]
  assign bb_for_body124_io_Out_26_ready = binaryOp_add2941_io_enable_ready; // @[extracted_function_conv.scala 893:30]
  assign bb_for_body124_io_Out_27_ready = Gep_arrayidx3042_io_enable_ready; // @[extracted_function_conv.scala 896:30]
  assign bb_for_body124_io_Out_28_ready = ld_43_io_enable_ready; // @[extracted_function_conv.scala 899:19]
  assign bb_for_body124_io_Out_29_ready = sextconv3244_io_enable_ready; // @[extracted_function_conv.scala 902:26]
  assign bb_for_body124_io_Out_30_ready = binaryOp_mul3345_io_enable_ready; // @[extracted_function_conv.scala 905:30]
  assign bb_for_body124_io_Out_31_ready = binaryOp_add3446_io_enable_ready; // @[extracted_function_conv.scala 908:30]
  assign bb_for_body124_io_Out_32_ready = st_47_io_enable_ready; // @[extracted_function_conv.scala 911:19]
  assign bb_for_body124_io_Out_33_ready = ld_48_io_enable_ready; // @[extracted_function_conv.scala 914:19]
  assign bb_for_body124_io_Out_34_ready = binaryOp_add4249_io_enable_ready; // @[extracted_function_conv.scala 917:30]
  assign bb_for_body124_io_Out_35_ready = Gep_arrayidx4350_io_enable_ready; // @[extracted_function_conv.scala 920:30]
  assign bb_for_body124_io_Out_36_ready = ld_51_io_enable_ready; // @[extracted_function_conv.scala 923:19]
  assign bb_for_body124_io_Out_37_ready = sextconv4552_io_enable_ready; // @[extracted_function_conv.scala 926:26]
  assign bb_for_body124_io_Out_38_ready = binaryOp_mul4653_io_enable_ready; // @[extracted_function_conv.scala 929:30]
  assign bb_for_body124_io_Out_39_ready = binaryOp_add4754_io_enable_ready; // @[extracted_function_conv.scala 932:30]
  assign bb_for_body124_io_Out_40_ready = st_55_io_enable_ready; // @[extracted_function_conv.scala 935:19]
  assign bb_for_body124_io_Out_41_ready = ld_56_io_enable_ready; // @[extracted_function_conv.scala 938:19]
  assign bb_for_body124_io_Out_42_ready = binaryOp_mul5257_io_enable_ready; // @[extracted_function_conv.scala 941:30]
  assign bb_for_body124_io_Out_43_ready = binaryOp_add5358_io_enable_ready; // @[extracted_function_conv.scala 944:30]
  assign bb_for_body124_io_Out_44_ready = Gep_arrayidx5459_io_enable_ready; // @[extracted_function_conv.scala 947:30]
  assign bb_for_body124_io_Out_45_ready = ld_60_io_enable_ready; // @[extracted_function_conv.scala 950:19]
  assign bb_for_body124_io_Out_46_ready = sextconv5661_io_enable_ready; // @[extracted_function_conv.scala 953:26]
  assign bb_for_body124_io_Out_47_ready = binaryOp_mul5762_io_enable_ready; // @[extracted_function_conv.scala 956:30]
  assign bb_for_body124_io_Out_48_ready = binaryOp_add5863_io_enable_ready; // @[extracted_function_conv.scala 959:30]
  assign bb_for_body124_io_Out_49_ready = st_64_io_enable_ready; // @[extracted_function_conv.scala 962:19]
  assign bb_for_body124_io_Out_50_ready = ld_65_io_enable_ready; // @[extracted_function_conv.scala 965:19]
  assign bb_for_body124_io_Out_51_ready = binaryOp_add6566_io_enable_ready; // @[extracted_function_conv.scala 968:30]
  assign bb_for_body124_io_Out_52_ready = Gep_arrayidx6667_io_enable_ready; // @[extracted_function_conv.scala 971:30]
  assign bb_for_body124_io_Out_53_ready = ld_68_io_enable_ready; // @[extracted_function_conv.scala 974:19]
  assign bb_for_body124_io_Out_54_ready = sextconv6869_io_enable_ready; // @[extracted_function_conv.scala 977:26]
  assign bb_for_body124_io_Out_55_ready = binaryOp_mul6970_io_enable_ready; // @[extracted_function_conv.scala 980:30]
  assign bb_for_body124_io_Out_56_ready = binaryOp_add7071_io_enable_ready; // @[extracted_function_conv.scala 983:30]
  assign bb_for_body124_io_Out_57_ready = st_72_io_enable_ready; // @[extracted_function_conv.scala 986:19]
  assign bb_for_body124_io_Out_58_ready = ld_73_io_enable_ready; // @[extracted_function_conv.scala 989:19]
  assign bb_for_body124_io_Out_59_ready = binaryOp_add7774_io_enable_ready; // @[extracted_function_conv.scala 992:30]
  assign bb_for_body124_io_Out_60_ready = Gep_arrayidx7875_io_enable_ready; // @[extracted_function_conv.scala 995:30]
  assign bb_for_body124_io_Out_61_ready = ld_76_io_enable_ready; // @[extracted_function_conv.scala 998:19]
  assign bb_for_body124_io_Out_62_ready = sextconv8077_io_enable_ready; // @[extracted_function_conv.scala 1001:26]
  assign bb_for_body124_io_Out_63_ready = binaryOp_mul8178_io_enable_ready; // @[extracted_function_conv.scala 1004:30]
  assign bb_for_body124_io_Out_64_ready = binaryOp_add8279_io_enable_ready; // @[extracted_function_conv.scala 1007:30]
  assign bb_for_body124_io_Out_65_ready = st_80_io_enable_ready; // @[extracted_function_conv.scala 1010:19]
  assign bb_for_body124_io_Out_66_ready = ld_81_io_enable_ready; // @[extracted_function_conv.scala 1013:19]
  assign bb_for_body124_io_Out_67_ready = binaryOp_add8882_io_enable_ready; // @[extracted_function_conv.scala 1016:30]
  assign bb_for_body124_io_Out_68_ready = Gep_arrayidx8983_io_enable_ready; // @[extracted_function_conv.scala 1019:30]
  assign bb_for_body124_io_Out_69_ready = ld_84_io_enable_ready; // @[extracted_function_conv.scala 1022:19]
  assign bb_for_body124_io_Out_70_ready = sextconv9185_io_enable_ready; // @[extracted_function_conv.scala 1025:26]
  assign bb_for_body124_io_Out_71_ready = binaryOp_mul9286_io_enable_ready; // @[extracted_function_conv.scala 1028:30]
  assign bb_for_body124_io_Out_72_ready = binaryOp_add9387_io_enable_ready; // @[extracted_function_conv.scala 1031:30]
  assign bb_for_body124_io_Out_73_ready = st_88_io_enable_ready; // @[extracted_function_conv.scala 1034:19]
  assign bb_for_body124_io_Out_74_ready = ld_89_io_enable_ready; // @[extracted_function_conv.scala 1037:19]
  assign bb_for_body124_io_Out_75_ready = binaryOp_add10090_io_enable_ready; // @[extracted_function_conv.scala 1040:31]
  assign bb_for_body124_io_Out_76_ready = Gep_arrayidx10191_io_enable_ready; // @[extracted_function_conv.scala 1043:31]
  assign bb_for_body124_io_Out_77_ready = ld_92_io_enable_ready; // @[extracted_function_conv.scala 1046:19]
  assign bb_for_body124_io_Out_78_ready = sextconv10393_io_enable_ready; // @[extracted_function_conv.scala 1049:27]
  assign bb_for_body124_io_Out_79_ready = binaryOp_mul10494_io_enable_ready; // @[extracted_function_conv.scala 1052:31]
  assign bb_for_body124_io_Out_80_ready = binaryOp_add10595_io_enable_ready; // @[extracted_function_conv.scala 1055:31]
  assign bb_for_body124_io_Out_81_ready = st_96_io_enable_ready; // @[extracted_function_conv.scala 1058:19]
  assign bb_for_body124_io_Out_82_ready = ld_97_io_enable_ready; // @[extracted_function_conv.scala 1061:19]
  assign bb_for_body124_io_Out_83_ready = binaryOp_add11298_io_enable_ready; // @[extracted_function_conv.scala 1064:31]
  assign bb_for_body124_io_Out_84_ready = Gep_arrayidx11399_io_enable_ready; // @[extracted_function_conv.scala 1067:31]
  assign bb_for_body124_io_Out_85_ready = ld_100_io_enable_ready; // @[extracted_function_conv.scala 1070:20]
  assign bb_for_body124_io_Out_86_ready = sextconv115101_io_enable_ready; // @[extracted_function_conv.scala 1073:28]
  assign bb_for_body124_io_Out_87_ready = binaryOp_mul116102_io_enable_ready; // @[extracted_function_conv.scala 1076:32]
  assign bb_for_body124_io_Out_88_ready = binaryOp_add117103_io_enable_ready; // @[extracted_function_conv.scala 1079:32]
  assign bb_for_body124_io_Out_89_ready = st_104_io_enable_ready; // @[extracted_function_conv.scala 1082:20]
  assign bb_for_body124_io_Out_90_ready = binaryOp_inc105_io_enable_ready; // @[extracted_function_conv.scala 1085:29]
  assign bb_for_body124_io_Out_91_ready = icmp_exitcond106_io_enable_ready; // @[extracted_function_conv.scala 1088:30]
  assign bb_for_body124_io_Out_92_ready = br_107_io_enable_ready; // @[extracted_function_conv.scala 1091:20]
  assign bb_for_body124_io_predicateIn_0_valid = Loop_0_io_activate_loop_back_valid; // @[extracted_function_conv.scala 520:36]
  assign bb_for_body124_io_predicateIn_0_bits_taskID = Loop_0_io_activate_loop_back_bits_taskID; // @[extracted_function_conv.scala 520:36]
  assign bb_for_body124_io_predicateIn_0_bits_control = Loop_0_io_activate_loop_back_bits_control; // @[extracted_function_conv.scala 520:36]
  assign bb_for_body124_io_predicateIn_1_valid = Loop_0_io_activate_loop_start_valid; // @[extracted_function_conv.scala 518:36]
  assign bb_for_body124_io_predicateIn_1_bits_taskID = Loop_0_io_activate_loop_start_bits_taskID; // @[extracted_function_conv.scala 518:36]
  assign bb_for_body124_io_predicateIn_1_bits_control = Loop_0_io_activate_loop_start_bits_control; // @[extracted_function_conv.scala 518:36]
  assign binaryOp_mul0_clock = clock;
  assign binaryOp_mul0_reset = reset;
  assign binaryOp_mul0_io_enable_valid = bb_entry0_io_Out_8_valid; // @[extracted_function_conv.scala 734:27]
  assign binaryOp_mul0_io_enable_bits_taskID = bb_entry0_io_Out_8_bits_taskID; // @[extracted_function_conv.scala 734:27]
  assign binaryOp_mul0_io_enable_bits_control = bb_entry0_io_Out_8_bits_control; // @[extracted_function_conv.scala 734:27]
  assign binaryOp_mul0_io_Out_0_ready = binaryOp_add1_io_LeftIO_ready; // @[extracted_function_conv.scala 1292:27]
  assign binaryOp_mul0_io_LeftIO_valid = InputSplitter_io_Out_data_field5_1_valid; // @[extracted_function_conv.scala 1536:27]
  assign binaryOp_mul0_io_LeftIO_bits_data = InputSplitter_io_Out_data_field5_1_bits_data; // @[extracted_function_conv.scala 1536:27]
  assign binaryOp_mul0_io_RightIO_valid = InputSplitter_io_Out_data_field4_0_valid; // @[extracted_function_conv.scala 1534:28]
  assign binaryOp_mul0_io_RightIO_bits_data = InputSplitter_io_Out_data_field4_0_bits_data; // @[extracted_function_conv.scala 1534:28]
  assign binaryOp_add1_clock = clock;
  assign binaryOp_add1_reset = reset;
  assign binaryOp_add1_io_enable_valid = bb_entry0_io_Out_9_valid; // @[extracted_function_conv.scala 737:27]
  assign binaryOp_add1_io_enable_bits_taskID = bb_entry0_io_Out_9_bits_taskID; // @[extracted_function_conv.scala 737:27]
  assign binaryOp_add1_io_enable_bits_control = bb_entry0_io_Out_9_bits_control; // @[extracted_function_conv.scala 737:27]
  assign binaryOp_add1_io_Out_0_ready = Loop_1_io_InLiveIn_1_ready; // @[extracted_function_conv.scala 592:25]
  assign binaryOp_add1_io_LeftIO_valid = binaryOp_mul0_io_Out_0_valid; // @[extracted_function_conv.scala 1292:27]
  assign binaryOp_add1_io_LeftIO_bits_data = binaryOp_mul0_io_Out_0_bits_data; // @[extracted_function_conv.scala 1292:27]
  assign binaryOp_add1_io_RightIO_valid = InputSplitter_io_Out_data_field3_0_valid; // @[extracted_function_conv.scala 1532:28]
  assign binaryOp_add1_io_RightIO_bits_data = InputSplitter_io_Out_data_field3_0_bits_data; // @[extracted_function_conv.scala 1532:28]
  assign Gep_arrayidx252_clock = clock;
  assign Gep_arrayidx252_reset = reset;
  assign Gep_arrayidx252_io_enable_valid = bb_entry0_io_Out_10_valid; // @[extracted_function_conv.scala 740:29]
  assign Gep_arrayidx252_io_enable_bits_taskID = bb_entry0_io_Out_10_bits_taskID; // @[extracted_function_conv.scala 740:29]
  assign Gep_arrayidx252_io_enable_bits_control = bb_entry0_io_Out_10_bits_control; // @[extracted_function_conv.scala 740:29]
  assign Gep_arrayidx252_io_Out_0_ready = Loop_1_io_InLiveIn_5_ready; // @[extracted_function_conv.scala 600:25]
  assign Gep_arrayidx252_io_baseAddress_valid = InputSplitter_io_Out_data_field1_1_valid; // @[extracted_function_conv.scala 1516:34]
  assign Gep_arrayidx252_io_baseAddress_bits_taskID = InputSplitter_io_Out_data_field1_1_bits_taskID; // @[extracted_function_conv.scala 1516:34]
  assign Gep_arrayidx252_io_baseAddress_bits_data = InputSplitter_io_Out_data_field1_1_bits_data; // @[extracted_function_conv.scala 1516:34]
  assign Gep_arrayidx252_io_idx_0_valid = const0_io_Out_valid; // @[extracted_function_conv.scala 1240:29]
  assign Gep_arrayidx383_clock = clock;
  assign Gep_arrayidx383_reset = reset;
  assign Gep_arrayidx383_io_enable_valid = bb_entry0_io_Out_11_valid; // @[extracted_function_conv.scala 743:29]
  assign Gep_arrayidx383_io_enable_bits_taskID = bb_entry0_io_Out_11_bits_taskID; // @[extracted_function_conv.scala 743:29]
  assign Gep_arrayidx383_io_enable_bits_control = bb_entry0_io_Out_11_bits_control; // @[extracted_function_conv.scala 743:29]
  assign Gep_arrayidx383_io_Out_0_ready = Loop_1_io_InLiveIn_6_ready; // @[extracted_function_conv.scala 602:25]
  assign Gep_arrayidx383_io_baseAddress_valid = InputSplitter_io_Out_data_field1_2_valid; // @[extracted_function_conv.scala 1518:34]
  assign Gep_arrayidx383_io_baseAddress_bits_taskID = InputSplitter_io_Out_data_field1_2_bits_taskID; // @[extracted_function_conv.scala 1518:34]
  assign Gep_arrayidx383_io_baseAddress_bits_data = InputSplitter_io_Out_data_field1_2_bits_data; // @[extracted_function_conv.scala 1518:34]
  assign Gep_arrayidx383_io_idx_0_valid = const1_io_Out_valid; // @[extracted_function_conv.scala 1242:29]
  assign Gep_arrayidx514_clock = clock;
  assign Gep_arrayidx514_reset = reset;
  assign Gep_arrayidx514_io_enable_valid = bb_entry0_io_Out_12_valid; // @[extracted_function_conv.scala 746:29]
  assign Gep_arrayidx514_io_enable_bits_taskID = bb_entry0_io_Out_12_bits_taskID; // @[extracted_function_conv.scala 746:29]
  assign Gep_arrayidx514_io_enable_bits_control = bb_entry0_io_Out_12_bits_control; // @[extracted_function_conv.scala 746:29]
  assign Gep_arrayidx514_io_Out_0_ready = Loop_1_io_InLiveIn_7_ready; // @[extracted_function_conv.scala 604:25]
  assign Gep_arrayidx514_io_baseAddress_valid = InputSplitter_io_Out_data_field1_3_valid; // @[extracted_function_conv.scala 1520:34]
  assign Gep_arrayidx514_io_baseAddress_bits_taskID = InputSplitter_io_Out_data_field1_3_bits_taskID; // @[extracted_function_conv.scala 1520:34]
  assign Gep_arrayidx514_io_baseAddress_bits_data = InputSplitter_io_Out_data_field1_3_bits_data; // @[extracted_function_conv.scala 1520:34]
  assign Gep_arrayidx514_io_idx_0_valid = const2_io_Out_valid; // @[extracted_function_conv.scala 1244:29]
  assign Gep_arrayidx625_clock = clock;
  assign Gep_arrayidx625_reset = reset;
  assign Gep_arrayidx625_io_enable_valid = bb_entry0_io_Out_13_valid; // @[extracted_function_conv.scala 749:29]
  assign Gep_arrayidx625_io_enable_bits_taskID = bb_entry0_io_Out_13_bits_taskID; // @[extracted_function_conv.scala 749:29]
  assign Gep_arrayidx625_io_enable_bits_control = bb_entry0_io_Out_13_bits_control; // @[extracted_function_conv.scala 749:29]
  assign Gep_arrayidx625_io_Out_0_ready = Loop_1_io_InLiveIn_8_ready; // @[extracted_function_conv.scala 606:25]
  assign Gep_arrayidx625_io_baseAddress_valid = InputSplitter_io_Out_data_field1_4_valid; // @[extracted_function_conv.scala 1522:34]
  assign Gep_arrayidx625_io_baseAddress_bits_taskID = InputSplitter_io_Out_data_field1_4_bits_taskID; // @[extracted_function_conv.scala 1522:34]
  assign Gep_arrayidx625_io_baseAddress_bits_data = InputSplitter_io_Out_data_field1_4_bits_data; // @[extracted_function_conv.scala 1522:34]
  assign Gep_arrayidx625_io_idx_0_valid = const3_io_Out_valid; // @[extracted_function_conv.scala 1246:29]
  assign Gep_arrayidx746_clock = clock;
  assign Gep_arrayidx746_reset = reset;
  assign Gep_arrayidx746_io_enable_valid = bb_entry0_io_Out_14_valid; // @[extracted_function_conv.scala 752:29]
  assign Gep_arrayidx746_io_enable_bits_taskID = bb_entry0_io_Out_14_bits_taskID; // @[extracted_function_conv.scala 752:29]
  assign Gep_arrayidx746_io_enable_bits_control = bb_entry0_io_Out_14_bits_control; // @[extracted_function_conv.scala 752:29]
  assign Gep_arrayidx746_io_Out_0_ready = Loop_1_io_InLiveIn_9_ready; // @[extracted_function_conv.scala 608:25]
  assign Gep_arrayidx746_io_baseAddress_valid = InputSplitter_io_Out_data_field1_5_valid; // @[extracted_function_conv.scala 1524:34]
  assign Gep_arrayidx746_io_baseAddress_bits_taskID = InputSplitter_io_Out_data_field1_5_bits_taskID; // @[extracted_function_conv.scala 1524:34]
  assign Gep_arrayidx746_io_baseAddress_bits_data = InputSplitter_io_Out_data_field1_5_bits_data; // @[extracted_function_conv.scala 1524:34]
  assign Gep_arrayidx746_io_idx_0_valid = const4_io_Out_valid; // @[extracted_function_conv.scala 1248:29]
  assign Gep_arrayidx867_clock = clock;
  assign Gep_arrayidx867_reset = reset;
  assign Gep_arrayidx867_io_enable_valid = bb_entry0_io_Out_15_valid; // @[extracted_function_conv.scala 755:29]
  assign Gep_arrayidx867_io_enable_bits_taskID = bb_entry0_io_Out_15_bits_taskID; // @[extracted_function_conv.scala 755:29]
  assign Gep_arrayidx867_io_enable_bits_control = bb_entry0_io_Out_15_bits_control; // @[extracted_function_conv.scala 755:29]
  assign Gep_arrayidx867_io_Out_0_ready = Loop_1_io_InLiveIn_10_ready; // @[extracted_function_conv.scala 610:26]
  assign Gep_arrayidx867_io_baseAddress_valid = InputSplitter_io_Out_data_field1_6_valid; // @[extracted_function_conv.scala 1526:34]
  assign Gep_arrayidx867_io_baseAddress_bits_taskID = InputSplitter_io_Out_data_field1_6_bits_taskID; // @[extracted_function_conv.scala 1526:34]
  assign Gep_arrayidx867_io_baseAddress_bits_data = InputSplitter_io_Out_data_field1_6_bits_data; // @[extracted_function_conv.scala 1526:34]
  assign Gep_arrayidx867_io_idx_0_valid = const5_io_Out_valid; // @[extracted_function_conv.scala 1250:29]
  assign Gep_arrayidx978_clock = clock;
  assign Gep_arrayidx978_reset = reset;
  assign Gep_arrayidx978_io_enable_valid = bb_entry0_io_Out_16_valid; // @[extracted_function_conv.scala 758:29]
  assign Gep_arrayidx978_io_enable_bits_taskID = bb_entry0_io_Out_16_bits_taskID; // @[extracted_function_conv.scala 758:29]
  assign Gep_arrayidx978_io_enable_bits_control = bb_entry0_io_Out_16_bits_control; // @[extracted_function_conv.scala 758:29]
  assign Gep_arrayidx978_io_Out_0_ready = Loop_1_io_InLiveIn_11_ready; // @[extracted_function_conv.scala 612:26]
  assign Gep_arrayidx978_io_baseAddress_valid = InputSplitter_io_Out_data_field1_7_valid; // @[extracted_function_conv.scala 1528:34]
  assign Gep_arrayidx978_io_baseAddress_bits_taskID = InputSplitter_io_Out_data_field1_7_bits_taskID; // @[extracted_function_conv.scala 1528:34]
  assign Gep_arrayidx978_io_baseAddress_bits_data = InputSplitter_io_Out_data_field1_7_bits_data; // @[extracted_function_conv.scala 1528:34]
  assign Gep_arrayidx978_io_idx_0_valid = const6_io_Out_valid; // @[extracted_function_conv.scala 1252:29]
  assign Gep_arrayidx1099_clock = clock;
  assign Gep_arrayidx1099_reset = reset;
  assign Gep_arrayidx1099_io_enable_valid = bb_entry0_io_Out_17_valid; // @[extracted_function_conv.scala 761:30]
  assign Gep_arrayidx1099_io_enable_bits_taskID = bb_entry0_io_Out_17_bits_taskID; // @[extracted_function_conv.scala 761:30]
  assign Gep_arrayidx1099_io_enable_bits_control = bb_entry0_io_Out_17_bits_control; // @[extracted_function_conv.scala 761:30]
  assign Gep_arrayidx1099_io_Out_0_ready = Loop_1_io_InLiveIn_12_ready; // @[extracted_function_conv.scala 614:26]
  assign Gep_arrayidx1099_io_baseAddress_valid = InputSplitter_io_Out_data_field1_8_valid; // @[extracted_function_conv.scala 1530:35]
  assign Gep_arrayidx1099_io_baseAddress_bits_taskID = InputSplitter_io_Out_data_field1_8_bits_taskID; // @[extracted_function_conv.scala 1530:35]
  assign Gep_arrayidx1099_io_baseAddress_bits_data = InputSplitter_io_Out_data_field1_8_bits_data; // @[extracted_function_conv.scala 1530:35]
  assign Gep_arrayidx1099_io_idx_0_valid = const7_io_Out_valid; // @[extracted_function_conv.scala 1254:30]
  assign br_10_clock = clock;
  assign br_10_reset = reset;
  assign br_10_io_enable_valid = bb_entry0_io_Out_18_valid; // @[extracted_function_conv.scala 764:19]
  assign br_10_io_enable_bits_taskID = bb_entry0_io_Out_18_bits_taskID; // @[extracted_function_conv.scala 764:19]
  assign br_10_io_enable_bits_control = bb_entry0_io_Out_18_bits_control; // @[extracted_function_conv.scala 764:19]
  assign br_10_io_Out_0_ready = Loop_1_io_enable_ready; // @[extracted_function_conv.scala 540:20]
  assign ret_11_clock = clock;
  assign ret_11_reset = reset;
  assign ret_11_io_In_enable_valid = bb_for_cond_cleanup1_io_Out_0_valid; // @[extracted_function_conv.scala 767:23]
  assign ret_11_io_In_enable_bits_taskID = bb_for_cond_cleanup1_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 767:23]
  assign ret_11_io_In_enable_bits_control = bb_for_cond_cleanup1_io_Out_0_bits_control; // @[extracted_function_conv.scala 767:23]
  assign ret_11_io_Out_ready = io_out_ready; // @[extracted_function_conv.scala 1562:10]
  assign phi_conv_s1_y_031312_clock = clock;
  assign phi_conv_s1_y_031312_reset = reset;
  assign phi_conv_s1_y_031312_io_enable_valid = bb_for_body2_io_Out_5_valid; // @[extracted_function_conv.scala 780:34]
  assign phi_conv_s1_y_031312_io_enable_bits_control = bb_for_body2_io_Out_5_bits_control; // @[extracted_function_conv.scala 780:34]
  assign phi_conv_s1_y_031312_io_InData_0_valid = const8_io_Out_valid; // @[extracted_function_conv.scala 1256:37]
  assign phi_conv_s1_y_031312_io_InData_0_bits_taskID = const8_io_Out_bits_taskID; // @[extracted_function_conv.scala 1256:37]
  assign phi_conv_s1_y_031312_io_InData_1_valid = Loop_1_io_CarryDepenOut_field0_0_valid; // @[extracted_function_conv.scala 710:37]
  assign phi_conv_s1_y_031312_io_InData_1_bits_taskID = Loop_1_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_conv.scala 710:37]
  assign phi_conv_s1_y_031312_io_InData_1_bits_data = Loop_1_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_conv.scala 710:37]
  assign phi_conv_s1_y_031312_io_Mask_valid = bb_for_body2_io_MaskBB_0_valid; // @[extracted_function_conv.scala 1100:32]
  assign phi_conv_s1_y_031312_io_Mask_bits = bb_for_body2_io_MaskBB_0_bits; // @[extracted_function_conv.scala 1100:32]
  assign phi_conv_s1_y_031312_io_Out_0_ready = binaryOp_mul113_io_LeftIO_ready; // @[extracted_function_conv.scala 1294:29]
  assign phi_conv_s1_y_031312_io_Out_1_ready = binaryOp_mul720_io_LeftIO_ready; // @[extracted_function_conv.scala 1296:29]
  assign phi_conv_s1_y_031312_io_Out_2_ready = binaryOp_mul821_io_LeftIO_ready; // @[extracted_function_conv.scala 1298:29]
  assign phi_conv_s1_y_031312_io_Out_3_ready = binaryOp_inc12023_io_LeftIO_ready; // @[extracted_function_conv.scala 1300:31]
  assign binaryOp_mul113_clock = clock;
  assign binaryOp_mul113_reset = reset;
  assign binaryOp_mul113_io_enable_valid = bb_for_body2_io_Out_6_valid; // @[extracted_function_conv.scala 783:29]
  assign binaryOp_mul113_io_enable_bits_taskID = bb_for_body2_io_Out_6_bits_taskID; // @[extracted_function_conv.scala 783:29]
  assign binaryOp_mul113_io_enable_bits_control = bb_for_body2_io_Out_6_bits_control; // @[extracted_function_conv.scala 783:29]
  assign binaryOp_mul113_io_Out_0_ready = binaryOp_add214_io_LeftIO_ready; // @[extracted_function_conv.scala 1302:29]
  assign binaryOp_mul113_io_Out_1_ready = binaryOp_add417_io_LeftIO_ready; // @[extracted_function_conv.scala 1304:29]
  assign binaryOp_mul113_io_LeftIO_valid = phi_conv_s1_y_031312_io_Out_0_valid; // @[extracted_function_conv.scala 1294:29]
  assign binaryOp_mul113_io_LeftIO_bits_data = phi_conv_s1_y_031312_io_Out_0_bits_data; // @[extracted_function_conv.scala 1294:29]
  assign binaryOp_mul113_io_RightIO_valid = const9_io_Out_valid; // @[extracted_function_conv.scala 1258:30]
  assign binaryOp_add214_clock = clock;
  assign binaryOp_add214_reset = reset;
  assign binaryOp_add214_io_enable_valid = bb_for_body2_io_Out_7_valid; // @[extracted_function_conv.scala 786:29]
  assign binaryOp_add214_io_enable_bits_taskID = bb_for_body2_io_Out_7_bits_taskID; // @[extracted_function_conv.scala 786:29]
  assign binaryOp_add214_io_enable_bits_control = bb_for_body2_io_Out_7_bits_control; // @[extracted_function_conv.scala 786:29]
  assign binaryOp_add214_io_Out_0_ready = binaryOp_mul315_io_LeftIO_ready; // @[extracted_function_conv.scala 1306:29]
  assign binaryOp_add214_io_LeftIO_valid = binaryOp_mul113_io_Out_0_valid; // @[extracted_function_conv.scala 1302:29]
  assign binaryOp_add214_io_LeftIO_bits_data = binaryOp_mul113_io_Out_0_bits_data; // @[extracted_function_conv.scala 1302:29]
  assign binaryOp_add214_io_RightIO_valid = const10_io_Out_valid; // @[extracted_function_conv.scala 1260:30]
  assign binaryOp_mul315_clock = clock;
  assign binaryOp_mul315_reset = reset;
  assign binaryOp_mul315_io_enable_valid = bb_for_body2_io_Out_8_valid; // @[extracted_function_conv.scala 789:29]
  assign binaryOp_mul315_io_enable_bits_taskID = bb_for_body2_io_Out_8_bits_taskID; // @[extracted_function_conv.scala 789:29]
  assign binaryOp_mul315_io_enable_bits_control = bb_for_body2_io_Out_8_bits_control; // @[extracted_function_conv.scala 789:29]
  assign binaryOp_mul315_io_Out_0_ready = binaryOp_sub16_io_LeftIO_ready; // @[extracted_function_conv.scala 1308:28]
  assign binaryOp_mul315_io_LeftIO_valid = binaryOp_add214_io_Out_0_valid; // @[extracted_function_conv.scala 1306:29]
  assign binaryOp_mul315_io_LeftIO_bits_data = binaryOp_add214_io_Out_0_bits_data; // @[extracted_function_conv.scala 1306:29]
  assign binaryOp_mul315_io_RightIO_valid = Loop_1_io_OutLiveIn_field0_0_valid; // @[extracted_function_conv.scala 670:30]
  assign binaryOp_mul315_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_conv.scala 670:30]
  assign binaryOp_sub16_clock = clock;
  assign binaryOp_sub16_reset = reset;
  assign binaryOp_sub16_io_enable_valid = bb_for_body2_io_Out_9_valid; // @[extracted_function_conv.scala 792:28]
  assign binaryOp_sub16_io_enable_bits_taskID = bb_for_body2_io_Out_9_bits_taskID; // @[extracted_function_conv.scala 792:28]
  assign binaryOp_sub16_io_enable_bits_control = bb_for_body2_io_Out_9_bits_control; // @[extracted_function_conv.scala 792:28]
  assign binaryOp_sub16_io_Out_0_ready = Loop_0_io_InLiveIn_2_ready; // @[extracted_function_conv.scala 562:25]
  assign binaryOp_sub16_io_LeftIO_valid = binaryOp_mul315_io_Out_0_valid; // @[extracted_function_conv.scala 1308:28]
  assign binaryOp_sub16_io_LeftIO_bits_data = binaryOp_mul315_io_Out_0_bits_data; // @[extracted_function_conv.scala 1308:28]
  assign binaryOp_sub16_io_RightIO_valid = Loop_1_io_OutLiveIn_field1_1_valid; // @[extracted_function_conv.scala 676:29]
  assign binaryOp_sub16_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field1_1_bits_data; // @[extracted_function_conv.scala 676:29]
  assign binaryOp_add417_clock = clock;
  assign binaryOp_add417_reset = reset;
  assign binaryOp_add417_io_enable_valid = bb_for_body2_io_Out_10_valid; // @[extracted_function_conv.scala 795:29]
  assign binaryOp_add417_io_enable_bits_taskID = bb_for_body2_io_Out_10_bits_taskID; // @[extracted_function_conv.scala 795:29]
  assign binaryOp_add417_io_enable_bits_control = bb_for_body2_io_Out_10_bits_control; // @[extracted_function_conv.scala 795:29]
  assign binaryOp_add417_io_Out_0_ready = binaryOp_mul518_io_LeftIO_ready; // @[extracted_function_conv.scala 1310:29]
  assign binaryOp_add417_io_LeftIO_valid = binaryOp_mul113_io_Out_1_valid; // @[extracted_function_conv.scala 1304:29]
  assign binaryOp_add417_io_LeftIO_bits_data = binaryOp_mul113_io_Out_1_bits_data; // @[extracted_function_conv.scala 1304:29]
  assign binaryOp_add417_io_RightIO_valid = const11_io_Out_valid; // @[extracted_function_conv.scala 1262:30]
  assign binaryOp_mul518_clock = clock;
  assign binaryOp_mul518_reset = reset;
  assign binaryOp_mul518_io_enable_valid = bb_for_body2_io_Out_11_valid; // @[extracted_function_conv.scala 798:29]
  assign binaryOp_mul518_io_enable_bits_taskID = bb_for_body2_io_Out_11_bits_taskID; // @[extracted_function_conv.scala 798:29]
  assign binaryOp_mul518_io_enable_bits_control = bb_for_body2_io_Out_11_bits_control; // @[extracted_function_conv.scala 798:29]
  assign binaryOp_mul518_io_Out_0_ready = binaryOp_sub619_io_LeftIO_ready; // @[extracted_function_conv.scala 1312:29]
  assign binaryOp_mul518_io_LeftIO_valid = binaryOp_add417_io_Out_0_valid; // @[extracted_function_conv.scala 1310:29]
  assign binaryOp_mul518_io_LeftIO_bits_data = binaryOp_add417_io_Out_0_bits_data; // @[extracted_function_conv.scala 1310:29]
  assign binaryOp_mul518_io_RightIO_valid = Loop_1_io_OutLiveIn_field0_1_valid; // @[extracted_function_conv.scala 672:30]
  assign binaryOp_mul518_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field0_1_bits_data; // @[extracted_function_conv.scala 672:30]
  assign binaryOp_sub619_clock = clock;
  assign binaryOp_sub619_reset = reset;
  assign binaryOp_sub619_io_enable_valid = bb_for_body2_io_Out_12_valid; // @[extracted_function_conv.scala 801:29]
  assign binaryOp_sub619_io_enable_bits_taskID = bb_for_body2_io_Out_12_bits_taskID; // @[extracted_function_conv.scala 801:29]
  assign binaryOp_sub619_io_enable_bits_control = bb_for_body2_io_Out_12_bits_control; // @[extracted_function_conv.scala 801:29]
  assign binaryOp_sub619_io_Out_0_ready = Loop_0_io_InLiveIn_3_ready; // @[extracted_function_conv.scala 564:25]
  assign binaryOp_sub619_io_LeftIO_valid = binaryOp_mul518_io_Out_0_valid; // @[extracted_function_conv.scala 1312:29]
  assign binaryOp_sub619_io_LeftIO_bits_data = binaryOp_mul518_io_Out_0_bits_data; // @[extracted_function_conv.scala 1312:29]
  assign binaryOp_sub619_io_RightIO_valid = Loop_1_io_OutLiveIn_field1_2_valid; // @[extracted_function_conv.scala 678:30]
  assign binaryOp_sub619_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field1_2_bits_data; // @[extracted_function_conv.scala 678:30]
  assign binaryOp_mul720_clock = clock;
  assign binaryOp_mul720_reset = reset;
  assign binaryOp_mul720_io_enable_valid = bb_for_body2_io_Out_13_valid; // @[extracted_function_conv.scala 804:29]
  assign binaryOp_mul720_io_enable_bits_taskID = bb_for_body2_io_Out_13_bits_taskID; // @[extracted_function_conv.scala 804:29]
  assign binaryOp_mul720_io_enable_bits_control = bb_for_body2_io_Out_13_bits_control; // @[extracted_function_conv.scala 804:29]
  assign binaryOp_mul720_io_Out_0_ready = Loop_0_io_InLiveIn_1_ready; // @[extracted_function_conv.scala 560:25]
  assign binaryOp_mul720_io_LeftIO_valid = phi_conv_s1_y_031312_io_Out_1_valid; // @[extracted_function_conv.scala 1296:29]
  assign binaryOp_mul720_io_LeftIO_bits_data = phi_conv_s1_y_031312_io_Out_1_bits_data; // @[extracted_function_conv.scala 1296:29]
  assign binaryOp_mul720_io_RightIO_valid = Loop_1_io_OutLiveIn_field0_2_valid; // @[extracted_function_conv.scala 674:30]
  assign binaryOp_mul720_io_RightIO_bits_data = Loop_1_io_OutLiveIn_field0_2_bits_data; // @[extracted_function_conv.scala 674:30]
  assign binaryOp_mul821_clock = clock;
  assign binaryOp_mul821_reset = reset;
  assign binaryOp_mul821_io_enable_valid = bb_for_body2_io_Out_14_valid; // @[extracted_function_conv.scala 807:29]
  assign binaryOp_mul821_io_enable_bits_taskID = bb_for_body2_io_Out_14_bits_taskID; // @[extracted_function_conv.scala 807:29]
  assign binaryOp_mul821_io_enable_bits_control = bb_for_body2_io_Out_14_bits_control; // @[extracted_function_conv.scala 807:29]
  assign binaryOp_mul821_io_Out_0_ready = Loop_0_io_InLiveIn_0_ready; // @[extracted_function_conv.scala 558:25]
  assign binaryOp_mul821_io_LeftIO_valid = phi_conv_s1_y_031312_io_Out_2_valid; // @[extracted_function_conv.scala 1298:29]
  assign binaryOp_mul821_io_LeftIO_bits_data = phi_conv_s1_y_031312_io_Out_2_bits_data; // @[extracted_function_conv.scala 1298:29]
  assign binaryOp_mul821_io_RightIO_valid = const12_io_Out_valid; // @[extracted_function_conv.scala 1264:30]
  assign br_22_clock = clock;
  assign br_22_reset = reset;
  assign br_22_io_enable_valid = bb_for_body2_io_Out_15_valid; // @[extracted_function_conv.scala 810:19]
  assign br_22_io_enable_bits_taskID = bb_for_body2_io_Out_15_bits_taskID; // @[extracted_function_conv.scala 810:19]
  assign br_22_io_enable_bits_control = bb_for_body2_io_Out_15_bits_control; // @[extracted_function_conv.scala 810:19]
  assign br_22_io_Out_0_ready = Loop_0_io_enable_ready; // @[extracted_function_conv.scala 534:20]
  assign binaryOp_inc12023_clock = clock;
  assign binaryOp_inc12023_reset = reset;
  assign binaryOp_inc12023_io_enable_valid = bb_for_cond_cleanup113_io_Out_2_valid; // @[extracted_function_conv.scala 817:31]
  assign binaryOp_inc12023_io_enable_bits_taskID = bb_for_cond_cleanup113_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 817:31]
  assign binaryOp_inc12023_io_enable_bits_control = bb_for_cond_cleanup113_io_Out_2_bits_control; // @[extracted_function_conv.scala 817:31]
  assign binaryOp_inc12023_io_Out_0_ready = Loop_1_io_CarryDepenIn_0_ready; // @[extracted_function_conv.scala 700:29]
  assign binaryOp_inc12023_io_Out_1_ready = icmp_exitcond31424_io_LeftIO_ready; // @[extracted_function_conv.scala 1314:32]
  assign binaryOp_inc12023_io_LeftIO_valid = phi_conv_s1_y_031312_io_Out_3_valid; // @[extracted_function_conv.scala 1300:31]
  assign binaryOp_inc12023_io_LeftIO_bits_data = phi_conv_s1_y_031312_io_Out_3_bits_data; // @[extracted_function_conv.scala 1300:31]
  assign binaryOp_inc12023_io_RightIO_valid = const13_io_Out_valid; // @[extracted_function_conv.scala 1266:32]
  assign icmp_exitcond31424_clock = clock;
  assign icmp_exitcond31424_reset = reset;
  assign icmp_exitcond31424_io_enable_valid = bb_for_cond_cleanup113_io_Out_3_valid; // @[extracted_function_conv.scala 820:32]
  assign icmp_exitcond31424_io_enable_bits_taskID = bb_for_cond_cleanup113_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 820:32]
  assign icmp_exitcond31424_io_enable_bits_control = bb_for_cond_cleanup113_io_Out_3_bits_control; // @[extracted_function_conv.scala 820:32]
  assign icmp_exitcond31424_io_Out_0_ready = br_25_io_CmpIO_ready; // @[extracted_function_conv.scala 1316:18]
  assign icmp_exitcond31424_io_LeftIO_valid = binaryOp_inc12023_io_Out_1_valid; // @[extracted_function_conv.scala 1314:32]
  assign icmp_exitcond31424_io_LeftIO_bits_data = binaryOp_inc12023_io_Out_1_bits_data; // @[extracted_function_conv.scala 1314:32]
  assign icmp_exitcond31424_io_RightIO_valid = const14_io_Out_valid; // @[extracted_function_conv.scala 1268:33]
  assign br_25_clock = clock;
  assign br_25_reset = reset;
  assign br_25_io_enable_valid = bb_for_cond_cleanup113_io_Out_4_valid; // @[extracted_function_conv.scala 823:19]
  assign br_25_io_enable_bits_taskID = bb_for_cond_cleanup113_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 823:19]
  assign br_25_io_enable_bits_control = bb_for_cond_cleanup113_io_Out_4_bits_control; // @[extracted_function_conv.scala 823:19]
  assign br_25_io_CmpIO_valid = icmp_exitcond31424_io_Out_0_valid; // @[extracted_function_conv.scala 1316:18]
  assign br_25_io_CmpIO_bits_taskID = icmp_exitcond31424_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1316:18]
  assign br_25_io_CmpIO_bits_data = icmp_exitcond31424_io_Out_0_bits_data; // @[extracted_function_conv.scala 1316:18]
  assign br_25_io_TrueOutput_0_ready = Loop_1_io_loopFinish_0_ready; // @[extracted_function_conv.scala 544:27]
  assign br_25_io_FalseOutput_0_ready = Loop_1_io_loopBack_0_ready; // @[extracted_function_conv.scala 542:25]
  assign phi_conv_s1_x_031226_clock = clock;
  assign phi_conv_s1_x_031226_reset = reset;
  assign phi_conv_s1_x_031226_io_enable_valid = bb_for_body124_io_Out_11_valid; // @[extracted_function_conv.scala 848:34]
  assign phi_conv_s1_x_031226_io_enable_bits_control = bb_for_body124_io_Out_11_bits_control; // @[extracted_function_conv.scala 848:34]
  assign phi_conv_s1_x_031226_io_InData_0_valid = const15_io_Out_valid; // @[extracted_function_conv.scala 1270:37]
  assign phi_conv_s1_x_031226_io_InData_0_bits_taskID = const15_io_Out_bits_taskID; // @[extracted_function_conv.scala 1270:37]
  assign phi_conv_s1_x_031226_io_InData_1_valid = Loop_0_io_CarryDepenOut_field0_0_valid; // @[extracted_function_conv.scala 708:37]
  assign phi_conv_s1_x_031226_io_InData_1_bits_taskID = Loop_0_io_CarryDepenOut_field0_0_bits_taskID; // @[extracted_function_conv.scala 708:37]
  assign phi_conv_s1_x_031226_io_InData_1_bits_data = Loop_0_io_CarryDepenOut_field0_0_bits_data; // @[extracted_function_conv.scala 708:37]
  assign phi_conv_s1_x_031226_io_Mask_valid = bb_for_body124_io_MaskBB_0_valid; // @[extracted_function_conv.scala 1102:32]
  assign phi_conv_s1_x_031226_io_Mask_bits = bb_for_body124_io_MaskBB_0_bits; // @[extracted_function_conv.scala 1102:32]
  assign phi_conv_s1_x_031226_io_Out_0_ready = binaryOp_add1327_io_LeftIO_ready; // @[extracted_function_conv.scala 1318:30]
  assign phi_conv_s1_x_031226_io_Out_1_ready = binaryOp_add1531_io_LeftIO_ready; // @[extracted_function_conv.scala 1320:30]
  assign phi_conv_s1_x_031226_io_Out_2_ready = binaryOp_mul5257_io_LeftIO_ready; // @[extracted_function_conv.scala 1322:30]
  assign phi_conv_s1_x_031226_io_Out_3_ready = binaryOp_inc105_io_LeftIO_ready; // @[extracted_function_conv.scala 1324:29]
  assign binaryOp_add1327_clock = clock;
  assign binaryOp_add1327_reset = reset;
  assign binaryOp_add1327_io_enable_valid = bb_for_body124_io_Out_12_valid; // @[extracted_function_conv.scala 851:30]
  assign binaryOp_add1327_io_enable_bits_taskID = bb_for_body124_io_Out_12_bits_taskID; // @[extracted_function_conv.scala 851:30]
  assign binaryOp_add1327_io_enable_bits_control = bb_for_body124_io_Out_12_bits_control; // @[extracted_function_conv.scala 851:30]
  assign binaryOp_add1327_io_Out_0_ready = Gep_arrayidx28_io_idx_0_ready; // @[extracted_function_conv.scala 1326:28]
  assign binaryOp_add1327_io_LeftIO_valid = phi_conv_s1_x_031226_io_Out_0_valid; // @[extracted_function_conv.scala 1318:30]
  assign binaryOp_add1327_io_LeftIO_bits_data = phi_conv_s1_x_031226_io_Out_0_bits_data; // @[extracted_function_conv.scala 1318:30]
  assign binaryOp_add1327_io_RightIO_valid = Loop_0_io_OutLiveIn_field0_0_valid; // @[extracted_function_conv.scala 622:31]
  assign binaryOp_add1327_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field0_0_bits_data; // @[extracted_function_conv.scala 622:31]
  assign Gep_arrayidx28_clock = clock;
  assign Gep_arrayidx28_reset = reset;
  assign Gep_arrayidx28_io_enable_valid = bb_for_body124_io_Out_13_valid; // @[extracted_function_conv.scala 854:28]
  assign Gep_arrayidx28_io_enable_bits_taskID = bb_for_body124_io_Out_13_bits_taskID; // @[extracted_function_conv.scala 854:28]
  assign Gep_arrayidx28_io_enable_bits_control = bb_for_body124_io_Out_13_bits_control; // @[extracted_function_conv.scala 854:28]
  assign Gep_arrayidx28_io_Out_0_ready = ld_29_io_GepAddr_ready; // @[extracted_function_conv.scala 1328:20]
  assign Gep_arrayidx28_io_Out_1_ready = st_39_io_GepAddr_ready; // @[extracted_function_conv.scala 1330:20]
  assign Gep_arrayidx28_io_Out_2_ready = st_47_io_GepAddr_ready; // @[extracted_function_conv.scala 1332:20]
  assign Gep_arrayidx28_io_Out_3_ready = st_55_io_GepAddr_ready; // @[extracted_function_conv.scala 1334:20]
  assign Gep_arrayidx28_io_Out_4_ready = st_64_io_GepAddr_ready; // @[extracted_function_conv.scala 1336:20]
  assign Gep_arrayidx28_io_Out_5_ready = st_72_io_GepAddr_ready; // @[extracted_function_conv.scala 1338:20]
  assign Gep_arrayidx28_io_Out_6_ready = st_80_io_GepAddr_ready; // @[extracted_function_conv.scala 1340:20]
  assign Gep_arrayidx28_io_Out_7_ready = st_88_io_GepAddr_ready; // @[extracted_function_conv.scala 1342:20]
  assign Gep_arrayidx28_io_Out_8_ready = st_96_io_GepAddr_ready; // @[extracted_function_conv.scala 1344:20]
  assign Gep_arrayidx28_io_Out_9_ready = st_104_io_GepAddr_ready; // @[extracted_function_conv.scala 1346:21]
  assign Gep_arrayidx28_io_baseAddress_valid = Loop_0_io_OutLiveIn_field11_0_valid; // @[extracted_function_conv.scala 660:33]
  assign Gep_arrayidx28_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field11_0_bits_taskID; // @[extracted_function_conv.scala 660:33]
  assign Gep_arrayidx28_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field11_0_bits_data; // @[extracted_function_conv.scala 660:33]
  assign Gep_arrayidx28_io_idx_0_valid = binaryOp_add1327_io_Out_0_valid; // @[extracted_function_conv.scala 1326:28]
  assign Gep_arrayidx28_io_idx_0_bits_data = binaryOp_add1327_io_Out_0_bits_data; // @[extracted_function_conv.scala 1326:28]
  assign ld_29_clock = clock;
  assign ld_29_reset = reset;
  assign ld_29_io_enable_valid = bb_for_body124_io_Out_14_valid; // @[extracted_function_conv.scala 857:19]
  assign ld_29_io_enable_bits_taskID = bb_for_body124_io_Out_14_bits_taskID; // @[extracted_function_conv.scala 857:19]
  assign ld_29_io_enable_bits_control = bb_for_body124_io_Out_14_bits_control; // @[extracted_function_conv.scala 857:19]
  assign ld_29_io_Out_0_ready = binaryOp_add2138_io_RightIO_ready; // @[extracted_function_conv.scala 1348:31]
  assign ld_29_io_GepAddr_valid = Gep_arrayidx28_io_Out_0_valid; // @[extracted_function_conv.scala 1328:20]
  assign ld_29_io_GepAddr_bits_predicate = Gep_arrayidx28_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1328:20]
  assign ld_29_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1328:20]
  assign ld_29_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_0_bits_data; // @[extracted_function_conv.scala 1328:20]
  assign ld_29_io_memReq_ready = MemCtrl_io_ReadIn_0_ready; // @[extracted_function_conv.scala 1116:24]
  assign ld_29_io_memResp_valid = MemCtrl_io_ReadOut_0_valid; // @[extracted_function_conv.scala 1118:20]
  assign ld_29_io_memResp_data = MemCtrl_io_ReadOut_0_data; // @[extracted_function_conv.scala 1118:20]
  assign ld_30_clock = clock;
  assign ld_30_reset = reset;
  assign ld_30_io_enable_valid = bb_for_body124_io_Out_15_valid; // @[extracted_function_conv.scala 860:19]
  assign ld_30_io_enable_bits_taskID = bb_for_body124_io_Out_15_bits_taskID; // @[extracted_function_conv.scala 860:19]
  assign ld_30_io_enable_bits_control = bb_for_body124_io_Out_15_bits_control; // @[extracted_function_conv.scala 860:19]
  assign ld_30_io_Out_0_ready = binaryOp_mul2037_io_LeftIO_ready; // @[extracted_function_conv.scala 1350:30]
  assign ld_30_io_GepAddr_valid = Loop_0_io_OutLiveIn_field14_0_valid; // @[extracted_function_conv.scala 666:20]
  assign ld_30_io_GepAddr_bits_predicate = Loop_0_io_OutLiveIn_field14_0_bits_predicate; // @[extracted_function_conv.scala 666:20]
  assign ld_30_io_GepAddr_bits_taskID = Loop_0_io_OutLiveIn_field14_0_bits_taskID; // @[extracted_function_conv.scala 666:20]
  assign ld_30_io_GepAddr_bits_data = Loop_0_io_OutLiveIn_field14_0_bits_data; // @[extracted_function_conv.scala 666:20]
  assign ld_30_io_memReq_ready = MemCtrl_io_ReadIn_1_ready; // @[extracted_function_conv.scala 1120:24]
  assign ld_30_io_memResp_valid = MemCtrl_io_ReadOut_1_valid; // @[extracted_function_conv.scala 1122:20]
  assign ld_30_io_memResp_data = MemCtrl_io_ReadOut_1_data; // @[extracted_function_conv.scala 1122:20]
  assign binaryOp_add1531_clock = clock;
  assign binaryOp_add1531_reset = reset;
  assign binaryOp_add1531_io_enable_valid = bb_for_body124_io_Out_16_valid; // @[extracted_function_conv.scala 863:30]
  assign binaryOp_add1531_io_enable_bits_taskID = bb_for_body124_io_Out_16_bits_taskID; // @[extracted_function_conv.scala 863:30]
  assign binaryOp_add1531_io_enable_bits_control = bb_for_body124_io_Out_16_bits_control; // @[extracted_function_conv.scala 863:30]
  assign binaryOp_add1531_io_Out_0_ready = binaryOp_mul1632_io_LeftIO_ready; // @[extracted_function_conv.scala 1352:30]
  assign binaryOp_add1531_io_LeftIO_valid = phi_conv_s1_x_031226_io_Out_1_valid; // @[extracted_function_conv.scala 1320:30]
  assign binaryOp_add1531_io_LeftIO_bits_data = phi_conv_s1_x_031226_io_Out_1_bits_data; // @[extracted_function_conv.scala 1320:30]
  assign binaryOp_add1531_io_RightIO_valid = Loop_0_io_OutLiveIn_field1_0_valid; // @[extracted_function_conv.scala 624:31]
  assign binaryOp_add1531_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field1_0_bits_data; // @[extracted_function_conv.scala 624:31]
  assign binaryOp_mul1632_clock = clock;
  assign binaryOp_mul1632_reset = reset;
  assign binaryOp_mul1632_io_enable_valid = bb_for_body124_io_Out_17_valid; // @[extracted_function_conv.scala 866:30]
  assign binaryOp_mul1632_io_enable_bits_taskID = bb_for_body124_io_Out_17_bits_taskID; // @[extracted_function_conv.scala 866:30]
  assign binaryOp_mul1632_io_enable_bits_control = bb_for_body124_io_Out_17_bits_control; // @[extracted_function_conv.scala 866:30]
  assign binaryOp_mul1632_io_Out_0_ready = binaryOp_sub1733_io_LeftIO_ready; // @[extracted_function_conv.scala 1354:30]
  assign binaryOp_mul1632_io_LeftIO_valid = binaryOp_add1531_io_Out_0_valid; // @[extracted_function_conv.scala 1352:30]
  assign binaryOp_mul1632_io_LeftIO_bits_data = binaryOp_add1531_io_Out_0_bits_data; // @[extracted_function_conv.scala 1352:30]
  assign binaryOp_mul1632_io_RightIO_valid = const16_io_Out_valid; // @[extracted_function_conv.scala 1272:31]
  assign binaryOp_sub1733_clock = clock;
  assign binaryOp_sub1733_reset = reset;
  assign binaryOp_sub1733_io_enable_valid = bb_for_body124_io_Out_18_valid; // @[extracted_function_conv.scala 869:30]
  assign binaryOp_sub1733_io_enable_bits_taskID = bb_for_body124_io_Out_18_bits_taskID; // @[extracted_function_conv.scala 869:30]
  assign binaryOp_sub1733_io_enable_bits_control = bb_for_body124_io_Out_18_bits_control; // @[extracted_function_conv.scala 869:30]
  assign binaryOp_sub1733_io_Out_0_ready = Gep_arrayidx1834_io_idx_0_ready; // @[extracted_function_conv.scala 1356:30]
  assign binaryOp_sub1733_io_Out_1_ready = binaryOp_add2941_io_LeftIO_ready; // @[extracted_function_conv.scala 1358:30]
  assign binaryOp_sub1733_io_Out_2_ready = binaryOp_add4249_io_LeftIO_ready; // @[extracted_function_conv.scala 1360:30]
  assign binaryOp_sub1733_io_LeftIO_valid = binaryOp_mul1632_io_Out_0_valid; // @[extracted_function_conv.scala 1354:30]
  assign binaryOp_sub1733_io_LeftIO_bits_data = binaryOp_mul1632_io_Out_0_bits_data; // @[extracted_function_conv.scala 1354:30]
  assign binaryOp_sub1733_io_RightIO_valid = Loop_0_io_OutLiveIn_field5_0_valid; // @[extracted_function_conv.scala 632:31]
  assign binaryOp_sub1733_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field5_0_bits_data; // @[extracted_function_conv.scala 632:31]
  assign Gep_arrayidx1834_clock = clock;
  assign Gep_arrayidx1834_reset = reset;
  assign Gep_arrayidx1834_io_enable_valid = bb_for_body124_io_Out_19_valid; // @[extracted_function_conv.scala 872:30]
  assign Gep_arrayidx1834_io_enable_bits_taskID = bb_for_body124_io_Out_19_bits_taskID; // @[extracted_function_conv.scala 872:30]
  assign Gep_arrayidx1834_io_enable_bits_control = bb_for_body124_io_Out_19_bits_control; // @[extracted_function_conv.scala 872:30]
  assign Gep_arrayidx1834_io_Out_0_ready = ld_35_io_GepAddr_ready; // @[extracted_function_conv.scala 1362:20]
  assign Gep_arrayidx1834_io_baseAddress_valid = Loop_0_io_OutLiveIn_field10_0_valid; // @[extracted_function_conv.scala 642:35]
  assign Gep_arrayidx1834_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field10_0_bits_taskID; // @[extracted_function_conv.scala 642:35]
  assign Gep_arrayidx1834_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field10_0_bits_data; // @[extracted_function_conv.scala 642:35]
  assign Gep_arrayidx1834_io_idx_0_valid = binaryOp_sub1733_io_Out_0_valid; // @[extracted_function_conv.scala 1356:30]
  assign Gep_arrayidx1834_io_idx_0_bits_data = binaryOp_sub1733_io_Out_0_bits_data; // @[extracted_function_conv.scala 1356:30]
  assign ld_35_clock = clock;
  assign ld_35_reset = reset;
  assign ld_35_io_enable_valid = bb_for_body124_io_Out_20_valid; // @[extracted_function_conv.scala 875:19]
  assign ld_35_io_enable_bits_taskID = bb_for_body124_io_Out_20_bits_taskID; // @[extracted_function_conv.scala 875:19]
  assign ld_35_io_enable_bits_control = bb_for_body124_io_Out_20_bits_control; // @[extracted_function_conv.scala 875:19]
  assign ld_35_io_Out_0_ready = sextconv1936_io_Input_ready; // @[extracted_function_conv.scala 1364:25]
  assign ld_35_io_GepAddr_valid = Gep_arrayidx1834_io_Out_0_valid; // @[extracted_function_conv.scala 1362:20]
  assign ld_35_io_GepAddr_bits_predicate = Gep_arrayidx1834_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1362:20]
  assign ld_35_io_GepAddr_bits_taskID = Gep_arrayidx1834_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1362:20]
  assign ld_35_io_GepAddr_bits_data = Gep_arrayidx1834_io_Out_0_bits_data; // @[extracted_function_conv.scala 1362:20]
  assign ld_35_io_memReq_ready = MemCtrl_io_ReadIn_2_ready; // @[extracted_function_conv.scala 1124:24]
  assign ld_35_io_memResp_valid = MemCtrl_io_ReadOut_2_valid; // @[extracted_function_conv.scala 1126:20]
  assign ld_35_io_memResp_data = MemCtrl_io_ReadOut_2_data; // @[extracted_function_conv.scala 1126:20]
  assign sextconv1936_clock = clock;
  assign sextconv1936_reset = reset;
  assign sextconv1936_io_Input_valid = ld_35_io_Out_0_valid; // @[extracted_function_conv.scala 1364:25]
  assign sextconv1936_io_Input_bits_data = ld_35_io_Out_0_bits_data; // @[extracted_function_conv.scala 1364:25]
  assign sextconv1936_io_enable_valid = bb_for_body124_io_Out_21_valid; // @[extracted_function_conv.scala 878:26]
  assign sextconv1936_io_enable_bits_taskID = bb_for_body124_io_Out_21_bits_taskID; // @[extracted_function_conv.scala 878:26]
  assign sextconv1936_io_Out_0_ready = binaryOp_mul2037_io_RightIO_ready; // @[extracted_function_conv.scala 1366:31]
  assign binaryOp_mul2037_clock = clock;
  assign binaryOp_mul2037_reset = reset;
  assign binaryOp_mul2037_io_enable_valid = bb_for_body124_io_Out_22_valid; // @[extracted_function_conv.scala 881:30]
  assign binaryOp_mul2037_io_enable_bits_taskID = bb_for_body124_io_Out_22_bits_taskID; // @[extracted_function_conv.scala 881:30]
  assign binaryOp_mul2037_io_enable_bits_control = bb_for_body124_io_Out_22_bits_control; // @[extracted_function_conv.scala 881:30]
  assign binaryOp_mul2037_io_Out_0_ready = binaryOp_add2138_io_LeftIO_ready; // @[extracted_function_conv.scala 1368:30]
  assign binaryOp_mul2037_io_LeftIO_valid = ld_30_io_Out_0_valid; // @[extracted_function_conv.scala 1350:30]
  assign binaryOp_mul2037_io_LeftIO_bits_data = ld_30_io_Out_0_bits_data; // @[extracted_function_conv.scala 1350:30]
  assign binaryOp_mul2037_io_RightIO_valid = sextconv1936_io_Out_0_valid; // @[extracted_function_conv.scala 1366:31]
  assign binaryOp_mul2037_io_RightIO_bits_data = sextconv1936_io_Out_0_bits_data; // @[extracted_function_conv.scala 1366:31]
  assign binaryOp_add2138_clock = clock;
  assign binaryOp_add2138_reset = reset;
  assign binaryOp_add2138_io_enable_valid = bb_for_body124_io_Out_23_valid; // @[extracted_function_conv.scala 884:30]
  assign binaryOp_add2138_io_enable_bits_taskID = bb_for_body124_io_Out_23_bits_taskID; // @[extracted_function_conv.scala 884:30]
  assign binaryOp_add2138_io_enable_bits_control = bb_for_body124_io_Out_23_bits_control; // @[extracted_function_conv.scala 884:30]
  assign binaryOp_add2138_io_Out_0_ready = st_39_io_inData_ready; // @[extracted_function_conv.scala 1370:19]
  assign binaryOp_add2138_io_Out_1_ready = binaryOp_add3446_io_RightIO_ready; // @[extracted_function_conv.scala 1372:31]
  assign binaryOp_add2138_io_LeftIO_valid = binaryOp_mul2037_io_Out_0_valid; // @[extracted_function_conv.scala 1368:30]
  assign binaryOp_add2138_io_LeftIO_bits_data = binaryOp_mul2037_io_Out_0_bits_data; // @[extracted_function_conv.scala 1368:30]
  assign binaryOp_add2138_io_RightIO_valid = ld_29_io_Out_0_valid; // @[extracted_function_conv.scala 1348:31]
  assign binaryOp_add2138_io_RightIO_bits_data = ld_29_io_Out_0_bits_data; // @[extracted_function_conv.scala 1348:31]
  assign st_39_clock = clock;
  assign st_39_reset = reset;
  assign st_39_io_enable_valid = bb_for_body124_io_Out_24_valid; // @[extracted_function_conv.scala 887:19]
  assign st_39_io_enable_bits_taskID = bb_for_body124_io_Out_24_bits_taskID; // @[extracted_function_conv.scala 887:19]
  assign st_39_io_enable_bits_control = bb_for_body124_io_Out_24_bits_control; // @[extracted_function_conv.scala 887:19]
  assign st_39_io_GepAddr_valid = Gep_arrayidx28_io_Out_1_valid; // @[extracted_function_conv.scala 1330:20]
  assign st_39_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 1330:20]
  assign st_39_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_1_bits_data; // @[extracted_function_conv.scala 1330:20]
  assign st_39_io_inData_valid = binaryOp_add2138_io_Out_0_valid; // @[extracted_function_conv.scala 1370:19]
  assign st_39_io_inData_bits_taskID = binaryOp_add2138_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1370:19]
  assign st_39_io_inData_bits_data = binaryOp_add2138_io_Out_0_bits_data; // @[extracted_function_conv.scala 1370:19]
  assign st_39_io_memReq_ready = MemCtrl_io_WriteIn_0_ready; // @[extracted_function_conv.scala 1128:25]
  assign st_39_io_memResp_valid = MemCtrl_io_WriteOut_0_valid; // @[extracted_function_conv.scala 1130:20]
  assign ld_40_clock = clock;
  assign ld_40_reset = reset;
  assign ld_40_io_enable_valid = bb_for_body124_io_Out_25_valid; // @[extracted_function_conv.scala 890:19]
  assign ld_40_io_enable_bits_taskID = bb_for_body124_io_Out_25_bits_taskID; // @[extracted_function_conv.scala 890:19]
  assign ld_40_io_enable_bits_control = bb_for_body124_io_Out_25_bits_control; // @[extracted_function_conv.scala 890:19]
  assign ld_40_io_Out_0_ready = binaryOp_mul3345_io_LeftIO_ready; // @[extracted_function_conv.scala 1374:30]
  assign ld_40_io_GepAddr_valid = Loop_0_io_OutLiveIn_field15_0_valid; // @[extracted_function_conv.scala 668:20]
  assign ld_40_io_GepAddr_bits_predicate = Loop_0_io_OutLiveIn_field15_0_bits_predicate; // @[extracted_function_conv.scala 668:20]
  assign ld_40_io_GepAddr_bits_taskID = Loop_0_io_OutLiveIn_field15_0_bits_taskID; // @[extracted_function_conv.scala 668:20]
  assign ld_40_io_GepAddr_bits_data = Loop_0_io_OutLiveIn_field15_0_bits_data; // @[extracted_function_conv.scala 668:20]
  assign ld_40_io_memReq_ready = MemCtrl_io_ReadIn_3_ready; // @[extracted_function_conv.scala 1132:24]
  assign ld_40_io_memResp_valid = MemCtrl_io_ReadOut_3_valid; // @[extracted_function_conv.scala 1134:20]
  assign ld_40_io_memResp_data = MemCtrl_io_ReadOut_3_data; // @[extracted_function_conv.scala 1134:20]
  assign binaryOp_add2941_clock = clock;
  assign binaryOp_add2941_reset = reset;
  assign binaryOp_add2941_io_enable_valid = bb_for_body124_io_Out_26_valid; // @[extracted_function_conv.scala 893:30]
  assign binaryOp_add2941_io_enable_bits_taskID = bb_for_body124_io_Out_26_bits_taskID; // @[extracted_function_conv.scala 893:30]
  assign binaryOp_add2941_io_enable_bits_control = bb_for_body124_io_Out_26_bits_control; // @[extracted_function_conv.scala 893:30]
  assign binaryOp_add2941_io_Out_0_ready = Gep_arrayidx3042_io_idx_0_ready; // @[extracted_function_conv.scala 1376:30]
  assign binaryOp_add2941_io_LeftIO_valid = binaryOp_sub1733_io_Out_1_valid; // @[extracted_function_conv.scala 1358:30]
  assign binaryOp_add2941_io_LeftIO_bits_data = binaryOp_sub1733_io_Out_1_bits_data; // @[extracted_function_conv.scala 1358:30]
  assign binaryOp_add2941_io_RightIO_valid = const17_io_Out_valid; // @[extracted_function_conv.scala 1274:31]
  assign Gep_arrayidx3042_clock = clock;
  assign Gep_arrayidx3042_reset = reset;
  assign Gep_arrayidx3042_io_enable_valid = bb_for_body124_io_Out_27_valid; // @[extracted_function_conv.scala 896:30]
  assign Gep_arrayidx3042_io_enable_bits_taskID = bb_for_body124_io_Out_27_bits_taskID; // @[extracted_function_conv.scala 896:30]
  assign Gep_arrayidx3042_io_enable_bits_control = bb_for_body124_io_Out_27_bits_control; // @[extracted_function_conv.scala 896:30]
  assign Gep_arrayidx3042_io_Out_0_ready = ld_43_io_GepAddr_ready; // @[extracted_function_conv.scala 1378:20]
  assign Gep_arrayidx3042_io_baseAddress_valid = Loop_0_io_OutLiveIn_field10_1_valid; // @[extracted_function_conv.scala 644:35]
  assign Gep_arrayidx3042_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field10_1_bits_taskID; // @[extracted_function_conv.scala 644:35]
  assign Gep_arrayidx3042_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field10_1_bits_data; // @[extracted_function_conv.scala 644:35]
  assign Gep_arrayidx3042_io_idx_0_valid = binaryOp_add2941_io_Out_0_valid; // @[extracted_function_conv.scala 1376:30]
  assign Gep_arrayidx3042_io_idx_0_bits_data = binaryOp_add2941_io_Out_0_bits_data; // @[extracted_function_conv.scala 1376:30]
  assign ld_43_clock = clock;
  assign ld_43_reset = reset;
  assign ld_43_io_enable_valid = bb_for_body124_io_Out_28_valid; // @[extracted_function_conv.scala 899:19]
  assign ld_43_io_enable_bits_taskID = bb_for_body124_io_Out_28_bits_taskID; // @[extracted_function_conv.scala 899:19]
  assign ld_43_io_enable_bits_control = bb_for_body124_io_Out_28_bits_control; // @[extracted_function_conv.scala 899:19]
  assign ld_43_io_Out_0_ready = sextconv3244_io_Input_ready; // @[extracted_function_conv.scala 1380:25]
  assign ld_43_io_GepAddr_valid = Gep_arrayidx3042_io_Out_0_valid; // @[extracted_function_conv.scala 1378:20]
  assign ld_43_io_GepAddr_bits_predicate = Gep_arrayidx3042_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1378:20]
  assign ld_43_io_GepAddr_bits_taskID = Gep_arrayidx3042_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1378:20]
  assign ld_43_io_GepAddr_bits_data = Gep_arrayidx3042_io_Out_0_bits_data; // @[extracted_function_conv.scala 1378:20]
  assign ld_43_io_memReq_ready = MemCtrl_io_ReadIn_4_ready; // @[extracted_function_conv.scala 1136:24]
  assign ld_43_io_memResp_valid = MemCtrl_io_ReadOut_4_valid; // @[extracted_function_conv.scala 1138:20]
  assign ld_43_io_memResp_data = MemCtrl_io_ReadOut_4_data; // @[extracted_function_conv.scala 1138:20]
  assign sextconv3244_clock = clock;
  assign sextconv3244_reset = reset;
  assign sextconv3244_io_Input_valid = ld_43_io_Out_0_valid; // @[extracted_function_conv.scala 1380:25]
  assign sextconv3244_io_Input_bits_data = ld_43_io_Out_0_bits_data; // @[extracted_function_conv.scala 1380:25]
  assign sextconv3244_io_enable_valid = bb_for_body124_io_Out_29_valid; // @[extracted_function_conv.scala 902:26]
  assign sextconv3244_io_enable_bits_taskID = bb_for_body124_io_Out_29_bits_taskID; // @[extracted_function_conv.scala 902:26]
  assign sextconv3244_io_Out_0_ready = binaryOp_mul3345_io_RightIO_ready; // @[extracted_function_conv.scala 1382:31]
  assign binaryOp_mul3345_clock = clock;
  assign binaryOp_mul3345_reset = reset;
  assign binaryOp_mul3345_io_enable_valid = bb_for_body124_io_Out_30_valid; // @[extracted_function_conv.scala 905:30]
  assign binaryOp_mul3345_io_enable_bits_taskID = bb_for_body124_io_Out_30_bits_taskID; // @[extracted_function_conv.scala 905:30]
  assign binaryOp_mul3345_io_enable_bits_control = bb_for_body124_io_Out_30_bits_control; // @[extracted_function_conv.scala 905:30]
  assign binaryOp_mul3345_io_Out_0_ready = binaryOp_add3446_io_LeftIO_ready; // @[extracted_function_conv.scala 1384:30]
  assign binaryOp_mul3345_io_LeftIO_valid = ld_40_io_Out_0_valid; // @[extracted_function_conv.scala 1374:30]
  assign binaryOp_mul3345_io_LeftIO_bits_data = ld_40_io_Out_0_bits_data; // @[extracted_function_conv.scala 1374:30]
  assign binaryOp_mul3345_io_RightIO_valid = sextconv3244_io_Out_0_valid; // @[extracted_function_conv.scala 1382:31]
  assign binaryOp_mul3345_io_RightIO_bits_data = sextconv3244_io_Out_0_bits_data; // @[extracted_function_conv.scala 1382:31]
  assign binaryOp_add3446_clock = clock;
  assign binaryOp_add3446_reset = reset;
  assign binaryOp_add3446_io_enable_valid = bb_for_body124_io_Out_31_valid; // @[extracted_function_conv.scala 908:30]
  assign binaryOp_add3446_io_enable_bits_taskID = bb_for_body124_io_Out_31_bits_taskID; // @[extracted_function_conv.scala 908:30]
  assign binaryOp_add3446_io_enable_bits_control = bb_for_body124_io_Out_31_bits_control; // @[extracted_function_conv.scala 908:30]
  assign binaryOp_add3446_io_Out_0_ready = st_47_io_inData_ready; // @[extracted_function_conv.scala 1386:19]
  assign binaryOp_add3446_io_Out_1_ready = binaryOp_add4754_io_RightIO_ready; // @[extracted_function_conv.scala 1388:31]
  assign binaryOp_add3446_io_LeftIO_valid = binaryOp_mul3345_io_Out_0_valid; // @[extracted_function_conv.scala 1384:30]
  assign binaryOp_add3446_io_LeftIO_bits_data = binaryOp_mul3345_io_Out_0_bits_data; // @[extracted_function_conv.scala 1384:30]
  assign binaryOp_add3446_io_RightIO_valid = binaryOp_add2138_io_Out_1_valid; // @[extracted_function_conv.scala 1372:31]
  assign binaryOp_add3446_io_RightIO_bits_data = binaryOp_add2138_io_Out_1_bits_data; // @[extracted_function_conv.scala 1372:31]
  assign st_47_clock = clock;
  assign st_47_reset = reset;
  assign st_47_io_enable_valid = bb_for_body124_io_Out_32_valid; // @[extracted_function_conv.scala 911:19]
  assign st_47_io_enable_bits_taskID = bb_for_body124_io_Out_32_bits_taskID; // @[extracted_function_conv.scala 911:19]
  assign st_47_io_enable_bits_control = bb_for_body124_io_Out_32_bits_control; // @[extracted_function_conv.scala 911:19]
  assign st_47_io_GepAddr_valid = Gep_arrayidx28_io_Out_2_valid; // @[extracted_function_conv.scala 1332:20]
  assign st_47_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 1332:20]
  assign st_47_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_2_bits_data; // @[extracted_function_conv.scala 1332:20]
  assign st_47_io_inData_valid = binaryOp_add3446_io_Out_0_valid; // @[extracted_function_conv.scala 1386:19]
  assign st_47_io_inData_bits_taskID = binaryOp_add3446_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1386:19]
  assign st_47_io_inData_bits_data = binaryOp_add3446_io_Out_0_bits_data; // @[extracted_function_conv.scala 1386:19]
  assign st_47_io_memReq_ready = MemCtrl_io_WriteIn_1_ready; // @[extracted_function_conv.scala 1140:25]
  assign st_47_io_memResp_valid = MemCtrl_io_WriteOut_1_valid; // @[extracted_function_conv.scala 1142:20]
  assign ld_48_clock = clock;
  assign ld_48_reset = reset;
  assign ld_48_io_enable_valid = bb_for_body124_io_Out_33_valid; // @[extracted_function_conv.scala 914:19]
  assign ld_48_io_enable_bits_taskID = bb_for_body124_io_Out_33_bits_taskID; // @[extracted_function_conv.scala 914:19]
  assign ld_48_io_enable_bits_control = bb_for_body124_io_Out_33_bits_control; // @[extracted_function_conv.scala 914:19]
  assign ld_48_io_Out_0_ready = binaryOp_mul4653_io_LeftIO_ready; // @[extracted_function_conv.scala 1390:30]
  assign ld_48_io_GepAddr_valid = Loop_0_io_OutLiveIn_field12_0_valid; // @[extracted_function_conv.scala 662:20]
  assign ld_48_io_GepAddr_bits_predicate = Loop_0_io_OutLiveIn_field12_0_bits_predicate; // @[extracted_function_conv.scala 662:20]
  assign ld_48_io_GepAddr_bits_taskID = Loop_0_io_OutLiveIn_field12_0_bits_taskID; // @[extracted_function_conv.scala 662:20]
  assign ld_48_io_GepAddr_bits_data = Loop_0_io_OutLiveIn_field12_0_bits_data; // @[extracted_function_conv.scala 662:20]
  assign ld_48_io_memReq_ready = MemCtrl_io_ReadIn_5_ready; // @[extracted_function_conv.scala 1144:24]
  assign ld_48_io_memResp_valid = MemCtrl_io_ReadOut_5_valid; // @[extracted_function_conv.scala 1146:20]
  assign ld_48_io_memResp_data = MemCtrl_io_ReadOut_5_data; // @[extracted_function_conv.scala 1146:20]
  assign binaryOp_add4249_clock = clock;
  assign binaryOp_add4249_reset = reset;
  assign binaryOp_add4249_io_enable_valid = bb_for_body124_io_Out_34_valid; // @[extracted_function_conv.scala 917:30]
  assign binaryOp_add4249_io_enable_bits_taskID = bb_for_body124_io_Out_34_bits_taskID; // @[extracted_function_conv.scala 917:30]
  assign binaryOp_add4249_io_enable_bits_control = bb_for_body124_io_Out_34_bits_control; // @[extracted_function_conv.scala 917:30]
  assign binaryOp_add4249_io_Out_0_ready = Gep_arrayidx4350_io_idx_0_ready; // @[extracted_function_conv.scala 1392:30]
  assign binaryOp_add4249_io_LeftIO_valid = binaryOp_sub1733_io_Out_2_valid; // @[extracted_function_conv.scala 1360:30]
  assign binaryOp_add4249_io_LeftIO_bits_data = binaryOp_sub1733_io_Out_2_bits_data; // @[extracted_function_conv.scala 1360:30]
  assign binaryOp_add4249_io_RightIO_valid = const18_io_Out_valid; // @[extracted_function_conv.scala 1276:31]
  assign Gep_arrayidx4350_clock = clock;
  assign Gep_arrayidx4350_reset = reset;
  assign Gep_arrayidx4350_io_enable_valid = bb_for_body124_io_Out_35_valid; // @[extracted_function_conv.scala 920:30]
  assign Gep_arrayidx4350_io_enable_bits_taskID = bb_for_body124_io_Out_35_bits_taskID; // @[extracted_function_conv.scala 920:30]
  assign Gep_arrayidx4350_io_enable_bits_control = bb_for_body124_io_Out_35_bits_control; // @[extracted_function_conv.scala 920:30]
  assign Gep_arrayidx4350_io_Out_0_ready = ld_51_io_GepAddr_ready; // @[extracted_function_conv.scala 1394:20]
  assign Gep_arrayidx4350_io_baseAddress_valid = Loop_0_io_OutLiveIn_field10_2_valid; // @[extracted_function_conv.scala 646:35]
  assign Gep_arrayidx4350_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field10_2_bits_taskID; // @[extracted_function_conv.scala 646:35]
  assign Gep_arrayidx4350_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field10_2_bits_data; // @[extracted_function_conv.scala 646:35]
  assign Gep_arrayidx4350_io_idx_0_valid = binaryOp_add4249_io_Out_0_valid; // @[extracted_function_conv.scala 1392:30]
  assign Gep_arrayidx4350_io_idx_0_bits_data = binaryOp_add4249_io_Out_0_bits_data; // @[extracted_function_conv.scala 1392:30]
  assign ld_51_clock = clock;
  assign ld_51_reset = reset;
  assign ld_51_io_enable_valid = bb_for_body124_io_Out_36_valid; // @[extracted_function_conv.scala 923:19]
  assign ld_51_io_enable_bits_taskID = bb_for_body124_io_Out_36_bits_taskID; // @[extracted_function_conv.scala 923:19]
  assign ld_51_io_enable_bits_control = bb_for_body124_io_Out_36_bits_control; // @[extracted_function_conv.scala 923:19]
  assign ld_51_io_Out_0_ready = sextconv4552_io_Input_ready; // @[extracted_function_conv.scala 1396:25]
  assign ld_51_io_GepAddr_valid = Gep_arrayidx4350_io_Out_0_valid; // @[extracted_function_conv.scala 1394:20]
  assign ld_51_io_GepAddr_bits_predicate = Gep_arrayidx4350_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1394:20]
  assign ld_51_io_GepAddr_bits_taskID = Gep_arrayidx4350_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1394:20]
  assign ld_51_io_GepAddr_bits_data = Gep_arrayidx4350_io_Out_0_bits_data; // @[extracted_function_conv.scala 1394:20]
  assign ld_51_io_memReq_ready = MemCtrl_io_ReadIn_6_ready; // @[extracted_function_conv.scala 1148:24]
  assign ld_51_io_memResp_valid = MemCtrl_io_ReadOut_6_valid; // @[extracted_function_conv.scala 1150:20]
  assign ld_51_io_memResp_data = MemCtrl_io_ReadOut_6_data; // @[extracted_function_conv.scala 1150:20]
  assign sextconv4552_clock = clock;
  assign sextconv4552_reset = reset;
  assign sextconv4552_io_Input_valid = ld_51_io_Out_0_valid; // @[extracted_function_conv.scala 1396:25]
  assign sextconv4552_io_Input_bits_data = ld_51_io_Out_0_bits_data; // @[extracted_function_conv.scala 1396:25]
  assign sextconv4552_io_enable_valid = bb_for_body124_io_Out_37_valid; // @[extracted_function_conv.scala 926:26]
  assign sextconv4552_io_enable_bits_taskID = bb_for_body124_io_Out_37_bits_taskID; // @[extracted_function_conv.scala 926:26]
  assign sextconv4552_io_Out_0_ready = binaryOp_mul4653_io_RightIO_ready; // @[extracted_function_conv.scala 1398:31]
  assign binaryOp_mul4653_clock = clock;
  assign binaryOp_mul4653_reset = reset;
  assign binaryOp_mul4653_io_enable_valid = bb_for_body124_io_Out_38_valid; // @[extracted_function_conv.scala 929:30]
  assign binaryOp_mul4653_io_enable_bits_taskID = bb_for_body124_io_Out_38_bits_taskID; // @[extracted_function_conv.scala 929:30]
  assign binaryOp_mul4653_io_enable_bits_control = bb_for_body124_io_Out_38_bits_control; // @[extracted_function_conv.scala 929:30]
  assign binaryOp_mul4653_io_Out_0_ready = binaryOp_add4754_io_LeftIO_ready; // @[extracted_function_conv.scala 1400:30]
  assign binaryOp_mul4653_io_LeftIO_valid = ld_48_io_Out_0_valid; // @[extracted_function_conv.scala 1390:30]
  assign binaryOp_mul4653_io_LeftIO_bits_data = ld_48_io_Out_0_bits_data; // @[extracted_function_conv.scala 1390:30]
  assign binaryOp_mul4653_io_RightIO_valid = sextconv4552_io_Out_0_valid; // @[extracted_function_conv.scala 1398:31]
  assign binaryOp_mul4653_io_RightIO_bits_data = sextconv4552_io_Out_0_bits_data; // @[extracted_function_conv.scala 1398:31]
  assign binaryOp_add4754_clock = clock;
  assign binaryOp_add4754_reset = reset;
  assign binaryOp_add4754_io_enable_valid = bb_for_body124_io_Out_39_valid; // @[extracted_function_conv.scala 932:30]
  assign binaryOp_add4754_io_enable_bits_taskID = bb_for_body124_io_Out_39_bits_taskID; // @[extracted_function_conv.scala 932:30]
  assign binaryOp_add4754_io_enable_bits_control = bb_for_body124_io_Out_39_bits_control; // @[extracted_function_conv.scala 932:30]
  assign binaryOp_add4754_io_Out_0_ready = st_55_io_inData_ready; // @[extracted_function_conv.scala 1402:19]
  assign binaryOp_add4754_io_Out_1_ready = binaryOp_add5863_io_RightIO_ready; // @[extracted_function_conv.scala 1404:31]
  assign binaryOp_add4754_io_LeftIO_valid = binaryOp_mul4653_io_Out_0_valid; // @[extracted_function_conv.scala 1400:30]
  assign binaryOp_add4754_io_LeftIO_bits_data = binaryOp_mul4653_io_Out_0_bits_data; // @[extracted_function_conv.scala 1400:30]
  assign binaryOp_add4754_io_RightIO_valid = binaryOp_add3446_io_Out_1_valid; // @[extracted_function_conv.scala 1388:31]
  assign binaryOp_add4754_io_RightIO_bits_data = binaryOp_add3446_io_Out_1_bits_data; // @[extracted_function_conv.scala 1388:31]
  assign st_55_clock = clock;
  assign st_55_reset = reset;
  assign st_55_io_enable_valid = bb_for_body124_io_Out_40_valid; // @[extracted_function_conv.scala 935:19]
  assign st_55_io_enable_bits_taskID = bb_for_body124_io_Out_40_bits_taskID; // @[extracted_function_conv.scala 935:19]
  assign st_55_io_enable_bits_control = bb_for_body124_io_Out_40_bits_control; // @[extracted_function_conv.scala 935:19]
  assign st_55_io_GepAddr_valid = Gep_arrayidx28_io_Out_3_valid; // @[extracted_function_conv.scala 1334:20]
  assign st_55_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 1334:20]
  assign st_55_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_3_bits_data; // @[extracted_function_conv.scala 1334:20]
  assign st_55_io_inData_valid = binaryOp_add4754_io_Out_0_valid; // @[extracted_function_conv.scala 1402:19]
  assign st_55_io_inData_bits_taskID = binaryOp_add4754_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1402:19]
  assign st_55_io_inData_bits_data = binaryOp_add4754_io_Out_0_bits_data; // @[extracted_function_conv.scala 1402:19]
  assign st_55_io_memReq_ready = MemCtrl_io_WriteIn_2_ready; // @[extracted_function_conv.scala 1152:25]
  assign st_55_io_memResp_valid = MemCtrl_io_WriteOut_2_valid; // @[extracted_function_conv.scala 1154:20]
  assign ld_56_clock = clock;
  assign ld_56_reset = reset;
  assign ld_56_io_enable_valid = bb_for_body124_io_Out_41_valid; // @[extracted_function_conv.scala 938:19]
  assign ld_56_io_enable_bits_taskID = bb_for_body124_io_Out_41_bits_taskID; // @[extracted_function_conv.scala 938:19]
  assign ld_56_io_enable_bits_control = bb_for_body124_io_Out_41_bits_control; // @[extracted_function_conv.scala 938:19]
  assign ld_56_io_Out_0_ready = binaryOp_mul5762_io_LeftIO_ready; // @[extracted_function_conv.scala 1406:30]
  assign ld_56_io_GepAddr_valid = Loop_0_io_OutLiveIn_field8_0_valid; // @[extracted_function_conv.scala 638:20]
  assign ld_56_io_GepAddr_bits_predicate = Loop_0_io_OutLiveIn_field8_0_bits_predicate; // @[extracted_function_conv.scala 638:20]
  assign ld_56_io_GepAddr_bits_taskID = Loop_0_io_OutLiveIn_field8_0_bits_taskID; // @[extracted_function_conv.scala 638:20]
  assign ld_56_io_GepAddr_bits_data = Loop_0_io_OutLiveIn_field8_0_bits_data; // @[extracted_function_conv.scala 638:20]
  assign ld_56_io_memReq_ready = MemCtrl_io_ReadIn_7_ready; // @[extracted_function_conv.scala 1156:24]
  assign ld_56_io_memResp_valid = MemCtrl_io_ReadOut_7_valid; // @[extracted_function_conv.scala 1158:20]
  assign ld_56_io_memResp_data = MemCtrl_io_ReadOut_7_data; // @[extracted_function_conv.scala 1158:20]
  assign binaryOp_mul5257_clock = clock;
  assign binaryOp_mul5257_reset = reset;
  assign binaryOp_mul5257_io_enable_valid = bb_for_body124_io_Out_42_valid; // @[extracted_function_conv.scala 941:30]
  assign binaryOp_mul5257_io_enable_bits_taskID = bb_for_body124_io_Out_42_bits_taskID; // @[extracted_function_conv.scala 941:30]
  assign binaryOp_mul5257_io_enable_bits_control = bb_for_body124_io_Out_42_bits_control; // @[extracted_function_conv.scala 941:30]
  assign binaryOp_mul5257_io_Out_0_ready = binaryOp_add5358_io_LeftIO_ready; // @[extracted_function_conv.scala 1408:30]
  assign binaryOp_mul5257_io_Out_1_ready = binaryOp_add8882_io_LeftIO_ready; // @[extracted_function_conv.scala 1410:30]
  assign binaryOp_mul5257_io_LeftIO_valid = phi_conv_s1_x_031226_io_Out_2_valid; // @[extracted_function_conv.scala 1322:30]
  assign binaryOp_mul5257_io_LeftIO_bits_data = phi_conv_s1_x_031226_io_Out_2_bits_data; // @[extracted_function_conv.scala 1322:30]
  assign binaryOp_mul5257_io_RightIO_valid = const19_io_Out_valid; // @[extracted_function_conv.scala 1278:31]
  assign binaryOp_add5358_clock = clock;
  assign binaryOp_add5358_reset = reset;
  assign binaryOp_add5358_io_enable_valid = bb_for_body124_io_Out_43_valid; // @[extracted_function_conv.scala 944:30]
  assign binaryOp_add5358_io_enable_bits_taskID = bb_for_body124_io_Out_43_bits_taskID; // @[extracted_function_conv.scala 944:30]
  assign binaryOp_add5358_io_enable_bits_control = bb_for_body124_io_Out_43_bits_control; // @[extracted_function_conv.scala 944:30]
  assign binaryOp_add5358_io_Out_0_ready = Gep_arrayidx5459_io_idx_0_ready; // @[extracted_function_conv.scala 1412:30]
  assign binaryOp_add5358_io_Out_1_ready = binaryOp_add6566_io_LeftIO_ready; // @[extracted_function_conv.scala 1414:30]
  assign binaryOp_add5358_io_Out_2_ready = binaryOp_add7774_io_LeftIO_ready; // @[extracted_function_conv.scala 1416:30]
  assign binaryOp_add5358_io_LeftIO_valid = binaryOp_mul5257_io_Out_0_valid; // @[extracted_function_conv.scala 1408:30]
  assign binaryOp_add5358_io_LeftIO_bits_data = binaryOp_mul5257_io_Out_0_bits_data; // @[extracted_function_conv.scala 1408:30]
  assign binaryOp_add5358_io_RightIO_valid = Loop_0_io_OutLiveIn_field2_0_valid; // @[extracted_function_conv.scala 626:31]
  assign binaryOp_add5358_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field2_0_bits_data; // @[extracted_function_conv.scala 626:31]
  assign Gep_arrayidx5459_clock = clock;
  assign Gep_arrayidx5459_reset = reset;
  assign Gep_arrayidx5459_io_enable_valid = bb_for_body124_io_Out_44_valid; // @[extracted_function_conv.scala 947:30]
  assign Gep_arrayidx5459_io_enable_bits_taskID = bb_for_body124_io_Out_44_bits_taskID; // @[extracted_function_conv.scala 947:30]
  assign Gep_arrayidx5459_io_enable_bits_control = bb_for_body124_io_Out_44_bits_control; // @[extracted_function_conv.scala 947:30]
  assign Gep_arrayidx5459_io_Out_0_ready = ld_60_io_GepAddr_ready; // @[extracted_function_conv.scala 1418:20]
  assign Gep_arrayidx5459_io_baseAddress_valid = Loop_0_io_OutLiveIn_field10_3_valid; // @[extracted_function_conv.scala 648:35]
  assign Gep_arrayidx5459_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field10_3_bits_taskID; // @[extracted_function_conv.scala 648:35]
  assign Gep_arrayidx5459_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field10_3_bits_data; // @[extracted_function_conv.scala 648:35]
  assign Gep_arrayidx5459_io_idx_0_valid = binaryOp_add5358_io_Out_0_valid; // @[extracted_function_conv.scala 1412:30]
  assign Gep_arrayidx5459_io_idx_0_bits_data = binaryOp_add5358_io_Out_0_bits_data; // @[extracted_function_conv.scala 1412:30]
  assign ld_60_clock = clock;
  assign ld_60_reset = reset;
  assign ld_60_io_enable_valid = bb_for_body124_io_Out_45_valid; // @[extracted_function_conv.scala 950:19]
  assign ld_60_io_enable_bits_taskID = bb_for_body124_io_Out_45_bits_taskID; // @[extracted_function_conv.scala 950:19]
  assign ld_60_io_enable_bits_control = bb_for_body124_io_Out_45_bits_control; // @[extracted_function_conv.scala 950:19]
  assign ld_60_io_Out_0_ready = sextconv5661_io_Input_ready; // @[extracted_function_conv.scala 1420:25]
  assign ld_60_io_GepAddr_valid = Gep_arrayidx5459_io_Out_0_valid; // @[extracted_function_conv.scala 1418:20]
  assign ld_60_io_GepAddr_bits_predicate = Gep_arrayidx5459_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1418:20]
  assign ld_60_io_GepAddr_bits_taskID = Gep_arrayidx5459_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1418:20]
  assign ld_60_io_GepAddr_bits_data = Gep_arrayidx5459_io_Out_0_bits_data; // @[extracted_function_conv.scala 1418:20]
  assign ld_60_io_memReq_ready = MemCtrl_io_ReadIn_8_ready; // @[extracted_function_conv.scala 1160:24]
  assign ld_60_io_memResp_valid = MemCtrl_io_ReadOut_8_valid; // @[extracted_function_conv.scala 1162:20]
  assign ld_60_io_memResp_data = MemCtrl_io_ReadOut_8_data; // @[extracted_function_conv.scala 1162:20]
  assign sextconv5661_clock = clock;
  assign sextconv5661_reset = reset;
  assign sextconv5661_io_Input_valid = ld_60_io_Out_0_valid; // @[extracted_function_conv.scala 1420:25]
  assign sextconv5661_io_Input_bits_data = ld_60_io_Out_0_bits_data; // @[extracted_function_conv.scala 1420:25]
  assign sextconv5661_io_enable_valid = bb_for_body124_io_Out_46_valid; // @[extracted_function_conv.scala 953:26]
  assign sextconv5661_io_enable_bits_taskID = bb_for_body124_io_Out_46_bits_taskID; // @[extracted_function_conv.scala 953:26]
  assign sextconv5661_io_Out_0_ready = binaryOp_mul5762_io_RightIO_ready; // @[extracted_function_conv.scala 1422:31]
  assign binaryOp_mul5762_clock = clock;
  assign binaryOp_mul5762_reset = reset;
  assign binaryOp_mul5762_io_enable_valid = bb_for_body124_io_Out_47_valid; // @[extracted_function_conv.scala 956:30]
  assign binaryOp_mul5762_io_enable_bits_taskID = bb_for_body124_io_Out_47_bits_taskID; // @[extracted_function_conv.scala 956:30]
  assign binaryOp_mul5762_io_enable_bits_control = bb_for_body124_io_Out_47_bits_control; // @[extracted_function_conv.scala 956:30]
  assign binaryOp_mul5762_io_Out_0_ready = binaryOp_add5863_io_LeftIO_ready; // @[extracted_function_conv.scala 1424:30]
  assign binaryOp_mul5762_io_LeftIO_valid = ld_56_io_Out_0_valid; // @[extracted_function_conv.scala 1406:30]
  assign binaryOp_mul5762_io_LeftIO_bits_data = ld_56_io_Out_0_bits_data; // @[extracted_function_conv.scala 1406:30]
  assign binaryOp_mul5762_io_RightIO_valid = sextconv5661_io_Out_0_valid; // @[extracted_function_conv.scala 1422:31]
  assign binaryOp_mul5762_io_RightIO_bits_data = sextconv5661_io_Out_0_bits_data; // @[extracted_function_conv.scala 1422:31]
  assign binaryOp_add5863_clock = clock;
  assign binaryOp_add5863_reset = reset;
  assign binaryOp_add5863_io_enable_valid = bb_for_body124_io_Out_48_valid; // @[extracted_function_conv.scala 959:30]
  assign binaryOp_add5863_io_enable_bits_taskID = bb_for_body124_io_Out_48_bits_taskID; // @[extracted_function_conv.scala 959:30]
  assign binaryOp_add5863_io_enable_bits_control = bb_for_body124_io_Out_48_bits_control; // @[extracted_function_conv.scala 959:30]
  assign binaryOp_add5863_io_Out_0_ready = st_64_io_inData_ready; // @[extracted_function_conv.scala 1426:19]
  assign binaryOp_add5863_io_Out_1_ready = binaryOp_add7071_io_RightIO_ready; // @[extracted_function_conv.scala 1428:31]
  assign binaryOp_add5863_io_LeftIO_valid = binaryOp_mul5762_io_Out_0_valid; // @[extracted_function_conv.scala 1424:30]
  assign binaryOp_add5863_io_LeftIO_bits_data = binaryOp_mul5762_io_Out_0_bits_data; // @[extracted_function_conv.scala 1424:30]
  assign binaryOp_add5863_io_RightIO_valid = binaryOp_add4754_io_Out_1_valid; // @[extracted_function_conv.scala 1404:31]
  assign binaryOp_add5863_io_RightIO_bits_data = binaryOp_add4754_io_Out_1_bits_data; // @[extracted_function_conv.scala 1404:31]
  assign st_64_clock = clock;
  assign st_64_reset = reset;
  assign st_64_io_enable_valid = bb_for_body124_io_Out_49_valid; // @[extracted_function_conv.scala 962:19]
  assign st_64_io_enable_bits_taskID = bb_for_body124_io_Out_49_bits_taskID; // @[extracted_function_conv.scala 962:19]
  assign st_64_io_enable_bits_control = bb_for_body124_io_Out_49_bits_control; // @[extracted_function_conv.scala 962:19]
  assign st_64_io_GepAddr_valid = Gep_arrayidx28_io_Out_4_valid; // @[extracted_function_conv.scala 1336:20]
  assign st_64_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 1336:20]
  assign st_64_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_4_bits_data; // @[extracted_function_conv.scala 1336:20]
  assign st_64_io_inData_valid = binaryOp_add5863_io_Out_0_valid; // @[extracted_function_conv.scala 1426:19]
  assign st_64_io_inData_bits_taskID = binaryOp_add5863_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1426:19]
  assign st_64_io_inData_bits_data = binaryOp_add5863_io_Out_0_bits_data; // @[extracted_function_conv.scala 1426:19]
  assign st_64_io_memReq_ready = MemCtrl_io_WriteIn_3_ready; // @[extracted_function_conv.scala 1164:25]
  assign st_64_io_memResp_valid = MemCtrl_io_WriteOut_3_valid; // @[extracted_function_conv.scala 1166:20]
  assign ld_65_clock = clock;
  assign ld_65_reset = reset;
  assign ld_65_io_enable_valid = bb_for_body124_io_Out_50_valid; // @[extracted_function_conv.scala 965:19]
  assign ld_65_io_enable_bits_taskID = bb_for_body124_io_Out_50_bits_taskID; // @[extracted_function_conv.scala 965:19]
  assign ld_65_io_enable_bits_control = bb_for_body124_io_Out_50_bits_control; // @[extracted_function_conv.scala 965:19]
  assign ld_65_io_Out_0_ready = binaryOp_mul6970_io_LeftIO_ready; // @[extracted_function_conv.scala 1430:30]
  assign ld_65_io_GepAddr_valid = Loop_0_io_OutLiveIn_field7_0_valid; // @[extracted_function_conv.scala 636:20]
  assign ld_65_io_GepAddr_bits_predicate = Loop_0_io_OutLiveIn_field7_0_bits_predicate; // @[extracted_function_conv.scala 636:20]
  assign ld_65_io_GepAddr_bits_taskID = Loop_0_io_OutLiveIn_field7_0_bits_taskID; // @[extracted_function_conv.scala 636:20]
  assign ld_65_io_GepAddr_bits_data = Loop_0_io_OutLiveIn_field7_0_bits_data; // @[extracted_function_conv.scala 636:20]
  assign ld_65_io_memReq_ready = MemCtrl_io_ReadIn_9_ready; // @[extracted_function_conv.scala 1168:24]
  assign ld_65_io_memResp_valid = MemCtrl_io_ReadOut_9_valid; // @[extracted_function_conv.scala 1170:20]
  assign ld_65_io_memResp_data = MemCtrl_io_ReadOut_9_data; // @[extracted_function_conv.scala 1170:20]
  assign binaryOp_add6566_clock = clock;
  assign binaryOp_add6566_reset = reset;
  assign binaryOp_add6566_io_enable_valid = bb_for_body124_io_Out_51_valid; // @[extracted_function_conv.scala 968:30]
  assign binaryOp_add6566_io_enable_bits_taskID = bb_for_body124_io_Out_51_bits_taskID; // @[extracted_function_conv.scala 968:30]
  assign binaryOp_add6566_io_enable_bits_control = bb_for_body124_io_Out_51_bits_control; // @[extracted_function_conv.scala 968:30]
  assign binaryOp_add6566_io_Out_0_ready = Gep_arrayidx6667_io_idx_0_ready; // @[extracted_function_conv.scala 1432:30]
  assign binaryOp_add6566_io_LeftIO_valid = binaryOp_add5358_io_Out_1_valid; // @[extracted_function_conv.scala 1414:30]
  assign binaryOp_add6566_io_LeftIO_bits_data = binaryOp_add5358_io_Out_1_bits_data; // @[extracted_function_conv.scala 1414:30]
  assign binaryOp_add6566_io_RightIO_valid = const20_io_Out_valid; // @[extracted_function_conv.scala 1280:31]
  assign Gep_arrayidx6667_clock = clock;
  assign Gep_arrayidx6667_reset = reset;
  assign Gep_arrayidx6667_io_enable_valid = bb_for_body124_io_Out_52_valid; // @[extracted_function_conv.scala 971:30]
  assign Gep_arrayidx6667_io_enable_bits_taskID = bb_for_body124_io_Out_52_bits_taskID; // @[extracted_function_conv.scala 971:30]
  assign Gep_arrayidx6667_io_enable_bits_control = bb_for_body124_io_Out_52_bits_control; // @[extracted_function_conv.scala 971:30]
  assign Gep_arrayidx6667_io_Out_0_ready = ld_68_io_GepAddr_ready; // @[extracted_function_conv.scala 1434:20]
  assign Gep_arrayidx6667_io_baseAddress_valid = Loop_0_io_OutLiveIn_field10_4_valid; // @[extracted_function_conv.scala 650:35]
  assign Gep_arrayidx6667_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field10_4_bits_taskID; // @[extracted_function_conv.scala 650:35]
  assign Gep_arrayidx6667_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field10_4_bits_data; // @[extracted_function_conv.scala 650:35]
  assign Gep_arrayidx6667_io_idx_0_valid = binaryOp_add6566_io_Out_0_valid; // @[extracted_function_conv.scala 1432:30]
  assign Gep_arrayidx6667_io_idx_0_bits_data = binaryOp_add6566_io_Out_0_bits_data; // @[extracted_function_conv.scala 1432:30]
  assign ld_68_clock = clock;
  assign ld_68_reset = reset;
  assign ld_68_io_enable_valid = bb_for_body124_io_Out_53_valid; // @[extracted_function_conv.scala 974:19]
  assign ld_68_io_enable_bits_taskID = bb_for_body124_io_Out_53_bits_taskID; // @[extracted_function_conv.scala 974:19]
  assign ld_68_io_enable_bits_control = bb_for_body124_io_Out_53_bits_control; // @[extracted_function_conv.scala 974:19]
  assign ld_68_io_Out_0_ready = sextconv6869_io_Input_ready; // @[extracted_function_conv.scala 1436:25]
  assign ld_68_io_GepAddr_valid = Gep_arrayidx6667_io_Out_0_valid; // @[extracted_function_conv.scala 1434:20]
  assign ld_68_io_GepAddr_bits_predicate = Gep_arrayidx6667_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1434:20]
  assign ld_68_io_GepAddr_bits_taskID = Gep_arrayidx6667_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1434:20]
  assign ld_68_io_GepAddr_bits_data = Gep_arrayidx6667_io_Out_0_bits_data; // @[extracted_function_conv.scala 1434:20]
  assign ld_68_io_memReq_ready = MemCtrl_io_ReadIn_10_ready; // @[extracted_function_conv.scala 1172:25]
  assign ld_68_io_memResp_valid = MemCtrl_io_ReadOut_10_valid; // @[extracted_function_conv.scala 1174:20]
  assign ld_68_io_memResp_data = MemCtrl_io_ReadOut_10_data; // @[extracted_function_conv.scala 1174:20]
  assign sextconv6869_clock = clock;
  assign sextconv6869_reset = reset;
  assign sextconv6869_io_Input_valid = ld_68_io_Out_0_valid; // @[extracted_function_conv.scala 1436:25]
  assign sextconv6869_io_Input_bits_data = ld_68_io_Out_0_bits_data; // @[extracted_function_conv.scala 1436:25]
  assign sextconv6869_io_enable_valid = bb_for_body124_io_Out_54_valid; // @[extracted_function_conv.scala 977:26]
  assign sextconv6869_io_enable_bits_taskID = bb_for_body124_io_Out_54_bits_taskID; // @[extracted_function_conv.scala 977:26]
  assign sextconv6869_io_Out_0_ready = binaryOp_mul6970_io_RightIO_ready; // @[extracted_function_conv.scala 1438:31]
  assign binaryOp_mul6970_clock = clock;
  assign binaryOp_mul6970_reset = reset;
  assign binaryOp_mul6970_io_enable_valid = bb_for_body124_io_Out_55_valid; // @[extracted_function_conv.scala 980:30]
  assign binaryOp_mul6970_io_enable_bits_taskID = bb_for_body124_io_Out_55_bits_taskID; // @[extracted_function_conv.scala 980:30]
  assign binaryOp_mul6970_io_enable_bits_control = bb_for_body124_io_Out_55_bits_control; // @[extracted_function_conv.scala 980:30]
  assign binaryOp_mul6970_io_Out_0_ready = binaryOp_add7071_io_LeftIO_ready; // @[extracted_function_conv.scala 1440:30]
  assign binaryOp_mul6970_io_LeftIO_valid = ld_65_io_Out_0_valid; // @[extracted_function_conv.scala 1430:30]
  assign binaryOp_mul6970_io_LeftIO_bits_data = ld_65_io_Out_0_bits_data; // @[extracted_function_conv.scala 1430:30]
  assign binaryOp_mul6970_io_RightIO_valid = sextconv6869_io_Out_0_valid; // @[extracted_function_conv.scala 1438:31]
  assign binaryOp_mul6970_io_RightIO_bits_data = sextconv6869_io_Out_0_bits_data; // @[extracted_function_conv.scala 1438:31]
  assign binaryOp_add7071_clock = clock;
  assign binaryOp_add7071_reset = reset;
  assign binaryOp_add7071_io_enable_valid = bb_for_body124_io_Out_56_valid; // @[extracted_function_conv.scala 983:30]
  assign binaryOp_add7071_io_enable_bits_taskID = bb_for_body124_io_Out_56_bits_taskID; // @[extracted_function_conv.scala 983:30]
  assign binaryOp_add7071_io_enable_bits_control = bb_for_body124_io_Out_56_bits_control; // @[extracted_function_conv.scala 983:30]
  assign binaryOp_add7071_io_Out_0_ready = st_72_io_inData_ready; // @[extracted_function_conv.scala 1442:19]
  assign binaryOp_add7071_io_Out_1_ready = binaryOp_add8279_io_RightIO_ready; // @[extracted_function_conv.scala 1444:31]
  assign binaryOp_add7071_io_LeftIO_valid = binaryOp_mul6970_io_Out_0_valid; // @[extracted_function_conv.scala 1440:30]
  assign binaryOp_add7071_io_LeftIO_bits_data = binaryOp_mul6970_io_Out_0_bits_data; // @[extracted_function_conv.scala 1440:30]
  assign binaryOp_add7071_io_RightIO_valid = binaryOp_add5863_io_Out_1_valid; // @[extracted_function_conv.scala 1428:31]
  assign binaryOp_add7071_io_RightIO_bits_data = binaryOp_add5863_io_Out_1_bits_data; // @[extracted_function_conv.scala 1428:31]
  assign st_72_clock = clock;
  assign st_72_reset = reset;
  assign st_72_io_enable_valid = bb_for_body124_io_Out_57_valid; // @[extracted_function_conv.scala 986:19]
  assign st_72_io_enable_bits_taskID = bb_for_body124_io_Out_57_bits_taskID; // @[extracted_function_conv.scala 986:19]
  assign st_72_io_enable_bits_control = bb_for_body124_io_Out_57_bits_control; // @[extracted_function_conv.scala 986:19]
  assign st_72_io_GepAddr_valid = Gep_arrayidx28_io_Out_5_valid; // @[extracted_function_conv.scala 1338:20]
  assign st_72_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_5_bits_taskID; // @[extracted_function_conv.scala 1338:20]
  assign st_72_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_5_bits_data; // @[extracted_function_conv.scala 1338:20]
  assign st_72_io_inData_valid = binaryOp_add7071_io_Out_0_valid; // @[extracted_function_conv.scala 1442:19]
  assign st_72_io_inData_bits_taskID = binaryOp_add7071_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1442:19]
  assign st_72_io_inData_bits_data = binaryOp_add7071_io_Out_0_bits_data; // @[extracted_function_conv.scala 1442:19]
  assign st_72_io_memReq_ready = MemCtrl_io_WriteIn_4_ready; // @[extracted_function_conv.scala 1176:25]
  assign st_72_io_memResp_valid = MemCtrl_io_WriteOut_4_valid; // @[extracted_function_conv.scala 1178:20]
  assign ld_73_clock = clock;
  assign ld_73_reset = reset;
  assign ld_73_io_enable_valid = bb_for_body124_io_Out_58_valid; // @[extracted_function_conv.scala 989:19]
  assign ld_73_io_enable_bits_taskID = bb_for_body124_io_Out_58_bits_taskID; // @[extracted_function_conv.scala 989:19]
  assign ld_73_io_enable_bits_control = bb_for_body124_io_Out_58_bits_control; // @[extracted_function_conv.scala 989:19]
  assign ld_73_io_Out_0_ready = binaryOp_mul8178_io_LeftIO_ready; // @[extracted_function_conv.scala 1446:30]
  assign ld_73_io_GepAddr_valid = Loop_0_io_OutLiveIn_field6_0_valid; // @[extracted_function_conv.scala 634:20]
  assign ld_73_io_GepAddr_bits_predicate = Loop_0_io_OutLiveIn_field6_0_bits_predicate; // @[extracted_function_conv.scala 634:20]
  assign ld_73_io_GepAddr_bits_taskID = Loop_0_io_OutLiveIn_field6_0_bits_taskID; // @[extracted_function_conv.scala 634:20]
  assign ld_73_io_GepAddr_bits_data = Loop_0_io_OutLiveIn_field6_0_bits_data; // @[extracted_function_conv.scala 634:20]
  assign ld_73_io_memReq_ready = MemCtrl_io_ReadIn_11_ready; // @[extracted_function_conv.scala 1180:25]
  assign ld_73_io_memResp_valid = MemCtrl_io_ReadOut_11_valid; // @[extracted_function_conv.scala 1182:20]
  assign ld_73_io_memResp_data = MemCtrl_io_ReadOut_11_data; // @[extracted_function_conv.scala 1182:20]
  assign binaryOp_add7774_clock = clock;
  assign binaryOp_add7774_reset = reset;
  assign binaryOp_add7774_io_enable_valid = bb_for_body124_io_Out_59_valid; // @[extracted_function_conv.scala 992:30]
  assign binaryOp_add7774_io_enable_bits_taskID = bb_for_body124_io_Out_59_bits_taskID; // @[extracted_function_conv.scala 992:30]
  assign binaryOp_add7774_io_enable_bits_control = bb_for_body124_io_Out_59_bits_control; // @[extracted_function_conv.scala 992:30]
  assign binaryOp_add7774_io_Out_0_ready = Gep_arrayidx7875_io_idx_0_ready; // @[extracted_function_conv.scala 1448:30]
  assign binaryOp_add7774_io_LeftIO_valid = binaryOp_add5358_io_Out_2_valid; // @[extracted_function_conv.scala 1416:30]
  assign binaryOp_add7774_io_LeftIO_bits_data = binaryOp_add5358_io_Out_2_bits_data; // @[extracted_function_conv.scala 1416:30]
  assign binaryOp_add7774_io_RightIO_valid = const21_io_Out_valid; // @[extracted_function_conv.scala 1282:31]
  assign Gep_arrayidx7875_clock = clock;
  assign Gep_arrayidx7875_reset = reset;
  assign Gep_arrayidx7875_io_enable_valid = bb_for_body124_io_Out_60_valid; // @[extracted_function_conv.scala 995:30]
  assign Gep_arrayidx7875_io_enable_bits_taskID = bb_for_body124_io_Out_60_bits_taskID; // @[extracted_function_conv.scala 995:30]
  assign Gep_arrayidx7875_io_enable_bits_control = bb_for_body124_io_Out_60_bits_control; // @[extracted_function_conv.scala 995:30]
  assign Gep_arrayidx7875_io_Out_0_ready = ld_76_io_GepAddr_ready; // @[extracted_function_conv.scala 1450:20]
  assign Gep_arrayidx7875_io_baseAddress_valid = Loop_0_io_OutLiveIn_field10_5_valid; // @[extracted_function_conv.scala 652:35]
  assign Gep_arrayidx7875_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field10_5_bits_taskID; // @[extracted_function_conv.scala 652:35]
  assign Gep_arrayidx7875_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field10_5_bits_data; // @[extracted_function_conv.scala 652:35]
  assign Gep_arrayidx7875_io_idx_0_valid = binaryOp_add7774_io_Out_0_valid; // @[extracted_function_conv.scala 1448:30]
  assign Gep_arrayidx7875_io_idx_0_bits_data = binaryOp_add7774_io_Out_0_bits_data; // @[extracted_function_conv.scala 1448:30]
  assign ld_76_clock = clock;
  assign ld_76_reset = reset;
  assign ld_76_io_enable_valid = bb_for_body124_io_Out_61_valid; // @[extracted_function_conv.scala 998:19]
  assign ld_76_io_enable_bits_taskID = bb_for_body124_io_Out_61_bits_taskID; // @[extracted_function_conv.scala 998:19]
  assign ld_76_io_enable_bits_control = bb_for_body124_io_Out_61_bits_control; // @[extracted_function_conv.scala 998:19]
  assign ld_76_io_Out_0_ready = sextconv8077_io_Input_ready; // @[extracted_function_conv.scala 1452:25]
  assign ld_76_io_GepAddr_valid = Gep_arrayidx7875_io_Out_0_valid; // @[extracted_function_conv.scala 1450:20]
  assign ld_76_io_GepAddr_bits_predicate = Gep_arrayidx7875_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1450:20]
  assign ld_76_io_GepAddr_bits_taskID = Gep_arrayidx7875_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1450:20]
  assign ld_76_io_GepAddr_bits_data = Gep_arrayidx7875_io_Out_0_bits_data; // @[extracted_function_conv.scala 1450:20]
  assign ld_76_io_memReq_ready = MemCtrl_io_ReadIn_12_ready; // @[extracted_function_conv.scala 1184:25]
  assign ld_76_io_memResp_valid = MemCtrl_io_ReadOut_12_valid; // @[extracted_function_conv.scala 1186:20]
  assign ld_76_io_memResp_data = MemCtrl_io_ReadOut_12_data; // @[extracted_function_conv.scala 1186:20]
  assign sextconv8077_clock = clock;
  assign sextconv8077_reset = reset;
  assign sextconv8077_io_Input_valid = ld_76_io_Out_0_valid; // @[extracted_function_conv.scala 1452:25]
  assign sextconv8077_io_Input_bits_data = ld_76_io_Out_0_bits_data; // @[extracted_function_conv.scala 1452:25]
  assign sextconv8077_io_enable_valid = bb_for_body124_io_Out_62_valid; // @[extracted_function_conv.scala 1001:26]
  assign sextconv8077_io_enable_bits_taskID = bb_for_body124_io_Out_62_bits_taskID; // @[extracted_function_conv.scala 1001:26]
  assign sextconv8077_io_Out_0_ready = binaryOp_mul8178_io_RightIO_ready; // @[extracted_function_conv.scala 1454:31]
  assign binaryOp_mul8178_clock = clock;
  assign binaryOp_mul8178_reset = reset;
  assign binaryOp_mul8178_io_enable_valid = bb_for_body124_io_Out_63_valid; // @[extracted_function_conv.scala 1004:30]
  assign binaryOp_mul8178_io_enable_bits_taskID = bb_for_body124_io_Out_63_bits_taskID; // @[extracted_function_conv.scala 1004:30]
  assign binaryOp_mul8178_io_enable_bits_control = bb_for_body124_io_Out_63_bits_control; // @[extracted_function_conv.scala 1004:30]
  assign binaryOp_mul8178_io_Out_0_ready = binaryOp_add8279_io_LeftIO_ready; // @[extracted_function_conv.scala 1456:30]
  assign binaryOp_mul8178_io_LeftIO_valid = ld_73_io_Out_0_valid; // @[extracted_function_conv.scala 1446:30]
  assign binaryOp_mul8178_io_LeftIO_bits_data = ld_73_io_Out_0_bits_data; // @[extracted_function_conv.scala 1446:30]
  assign binaryOp_mul8178_io_RightIO_valid = sextconv8077_io_Out_0_valid; // @[extracted_function_conv.scala 1454:31]
  assign binaryOp_mul8178_io_RightIO_bits_data = sextconv8077_io_Out_0_bits_data; // @[extracted_function_conv.scala 1454:31]
  assign binaryOp_add8279_clock = clock;
  assign binaryOp_add8279_reset = reset;
  assign binaryOp_add8279_io_enable_valid = bb_for_body124_io_Out_64_valid; // @[extracted_function_conv.scala 1007:30]
  assign binaryOp_add8279_io_enable_bits_taskID = bb_for_body124_io_Out_64_bits_taskID; // @[extracted_function_conv.scala 1007:30]
  assign binaryOp_add8279_io_enable_bits_control = bb_for_body124_io_Out_64_bits_control; // @[extracted_function_conv.scala 1007:30]
  assign binaryOp_add8279_io_Out_0_ready = st_80_io_inData_ready; // @[extracted_function_conv.scala 1458:19]
  assign binaryOp_add8279_io_Out_1_ready = binaryOp_add9387_io_RightIO_ready; // @[extracted_function_conv.scala 1460:31]
  assign binaryOp_add8279_io_LeftIO_valid = binaryOp_mul8178_io_Out_0_valid; // @[extracted_function_conv.scala 1456:30]
  assign binaryOp_add8279_io_LeftIO_bits_data = binaryOp_mul8178_io_Out_0_bits_data; // @[extracted_function_conv.scala 1456:30]
  assign binaryOp_add8279_io_RightIO_valid = binaryOp_add7071_io_Out_1_valid; // @[extracted_function_conv.scala 1444:31]
  assign binaryOp_add8279_io_RightIO_bits_data = binaryOp_add7071_io_Out_1_bits_data; // @[extracted_function_conv.scala 1444:31]
  assign st_80_clock = clock;
  assign st_80_reset = reset;
  assign st_80_io_enable_valid = bb_for_body124_io_Out_65_valid; // @[extracted_function_conv.scala 1010:19]
  assign st_80_io_enable_bits_taskID = bb_for_body124_io_Out_65_bits_taskID; // @[extracted_function_conv.scala 1010:19]
  assign st_80_io_enable_bits_control = bb_for_body124_io_Out_65_bits_control; // @[extracted_function_conv.scala 1010:19]
  assign st_80_io_GepAddr_valid = Gep_arrayidx28_io_Out_6_valid; // @[extracted_function_conv.scala 1340:20]
  assign st_80_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_6_bits_taskID; // @[extracted_function_conv.scala 1340:20]
  assign st_80_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_6_bits_data; // @[extracted_function_conv.scala 1340:20]
  assign st_80_io_inData_valid = binaryOp_add8279_io_Out_0_valid; // @[extracted_function_conv.scala 1458:19]
  assign st_80_io_inData_bits_taskID = binaryOp_add8279_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1458:19]
  assign st_80_io_inData_bits_data = binaryOp_add8279_io_Out_0_bits_data; // @[extracted_function_conv.scala 1458:19]
  assign st_80_io_memReq_ready = MemCtrl_io_WriteIn_5_ready; // @[extracted_function_conv.scala 1188:25]
  assign st_80_io_memResp_valid = MemCtrl_io_WriteOut_5_valid; // @[extracted_function_conv.scala 1190:20]
  assign ld_81_clock = clock;
  assign ld_81_reset = reset;
  assign ld_81_io_enable_valid = bb_for_body124_io_Out_66_valid; // @[extracted_function_conv.scala 1013:19]
  assign ld_81_io_enable_bits_taskID = bb_for_body124_io_Out_66_bits_taskID; // @[extracted_function_conv.scala 1013:19]
  assign ld_81_io_enable_bits_control = bb_for_body124_io_Out_66_bits_control; // @[extracted_function_conv.scala 1013:19]
  assign ld_81_io_Out_0_ready = binaryOp_mul9286_io_LeftIO_ready; // @[extracted_function_conv.scala 1462:30]
  assign ld_81_io_GepAddr_valid = Loop_0_io_OutLiveIn_field13_0_valid; // @[extracted_function_conv.scala 664:20]
  assign ld_81_io_GepAddr_bits_predicate = Loop_0_io_OutLiveIn_field13_0_bits_predicate; // @[extracted_function_conv.scala 664:20]
  assign ld_81_io_GepAddr_bits_taskID = Loop_0_io_OutLiveIn_field13_0_bits_taskID; // @[extracted_function_conv.scala 664:20]
  assign ld_81_io_GepAddr_bits_data = Loop_0_io_OutLiveIn_field13_0_bits_data; // @[extracted_function_conv.scala 664:20]
  assign ld_81_io_memReq_ready = MemCtrl_io_ReadIn_13_ready; // @[extracted_function_conv.scala 1192:25]
  assign ld_81_io_memResp_valid = MemCtrl_io_ReadOut_13_valid; // @[extracted_function_conv.scala 1194:20]
  assign ld_81_io_memResp_data = MemCtrl_io_ReadOut_13_data; // @[extracted_function_conv.scala 1194:20]
  assign binaryOp_add8882_clock = clock;
  assign binaryOp_add8882_reset = reset;
  assign binaryOp_add8882_io_enable_valid = bb_for_body124_io_Out_67_valid; // @[extracted_function_conv.scala 1016:30]
  assign binaryOp_add8882_io_enable_bits_taskID = bb_for_body124_io_Out_67_bits_taskID; // @[extracted_function_conv.scala 1016:30]
  assign binaryOp_add8882_io_enable_bits_control = bb_for_body124_io_Out_67_bits_control; // @[extracted_function_conv.scala 1016:30]
  assign binaryOp_add8882_io_Out_0_ready = Gep_arrayidx8983_io_idx_0_ready; // @[extracted_function_conv.scala 1464:30]
  assign binaryOp_add8882_io_Out_1_ready = binaryOp_add10090_io_LeftIO_ready; // @[extracted_function_conv.scala 1466:31]
  assign binaryOp_add8882_io_Out_2_ready = binaryOp_add11298_io_LeftIO_ready; // @[extracted_function_conv.scala 1468:31]
  assign binaryOp_add8882_io_LeftIO_valid = binaryOp_mul5257_io_Out_1_valid; // @[extracted_function_conv.scala 1410:30]
  assign binaryOp_add8882_io_LeftIO_bits_data = binaryOp_mul5257_io_Out_1_bits_data; // @[extracted_function_conv.scala 1410:30]
  assign binaryOp_add8882_io_RightIO_valid = Loop_0_io_OutLiveIn_field3_0_valid; // @[extracted_function_conv.scala 628:31]
  assign binaryOp_add8882_io_RightIO_bits_data = Loop_0_io_OutLiveIn_field3_0_bits_data; // @[extracted_function_conv.scala 628:31]
  assign Gep_arrayidx8983_clock = clock;
  assign Gep_arrayidx8983_reset = reset;
  assign Gep_arrayidx8983_io_enable_valid = bb_for_body124_io_Out_68_valid; // @[extracted_function_conv.scala 1019:30]
  assign Gep_arrayidx8983_io_enable_bits_taskID = bb_for_body124_io_Out_68_bits_taskID; // @[extracted_function_conv.scala 1019:30]
  assign Gep_arrayidx8983_io_enable_bits_control = bb_for_body124_io_Out_68_bits_control; // @[extracted_function_conv.scala 1019:30]
  assign Gep_arrayidx8983_io_Out_0_ready = ld_84_io_GepAddr_ready; // @[extracted_function_conv.scala 1470:20]
  assign Gep_arrayidx8983_io_baseAddress_valid = Loop_0_io_OutLiveIn_field10_6_valid; // @[extracted_function_conv.scala 654:35]
  assign Gep_arrayidx8983_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field10_6_bits_taskID; // @[extracted_function_conv.scala 654:35]
  assign Gep_arrayidx8983_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field10_6_bits_data; // @[extracted_function_conv.scala 654:35]
  assign Gep_arrayidx8983_io_idx_0_valid = binaryOp_add8882_io_Out_0_valid; // @[extracted_function_conv.scala 1464:30]
  assign Gep_arrayidx8983_io_idx_0_bits_data = binaryOp_add8882_io_Out_0_bits_data; // @[extracted_function_conv.scala 1464:30]
  assign ld_84_clock = clock;
  assign ld_84_reset = reset;
  assign ld_84_io_enable_valid = bb_for_body124_io_Out_69_valid; // @[extracted_function_conv.scala 1022:19]
  assign ld_84_io_enable_bits_taskID = bb_for_body124_io_Out_69_bits_taskID; // @[extracted_function_conv.scala 1022:19]
  assign ld_84_io_enable_bits_control = bb_for_body124_io_Out_69_bits_control; // @[extracted_function_conv.scala 1022:19]
  assign ld_84_io_Out_0_ready = sextconv9185_io_Input_ready; // @[extracted_function_conv.scala 1472:25]
  assign ld_84_io_GepAddr_valid = Gep_arrayidx8983_io_Out_0_valid; // @[extracted_function_conv.scala 1470:20]
  assign ld_84_io_GepAddr_bits_predicate = Gep_arrayidx8983_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1470:20]
  assign ld_84_io_GepAddr_bits_taskID = Gep_arrayidx8983_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1470:20]
  assign ld_84_io_GepAddr_bits_data = Gep_arrayidx8983_io_Out_0_bits_data; // @[extracted_function_conv.scala 1470:20]
  assign ld_84_io_memReq_ready = MemCtrl_io_ReadIn_14_ready; // @[extracted_function_conv.scala 1196:25]
  assign ld_84_io_memResp_valid = MemCtrl_io_ReadOut_14_valid; // @[extracted_function_conv.scala 1198:20]
  assign ld_84_io_memResp_data = MemCtrl_io_ReadOut_14_data; // @[extracted_function_conv.scala 1198:20]
  assign sextconv9185_clock = clock;
  assign sextconv9185_reset = reset;
  assign sextconv9185_io_Input_valid = ld_84_io_Out_0_valid; // @[extracted_function_conv.scala 1472:25]
  assign sextconv9185_io_Input_bits_data = ld_84_io_Out_0_bits_data; // @[extracted_function_conv.scala 1472:25]
  assign sextconv9185_io_enable_valid = bb_for_body124_io_Out_70_valid; // @[extracted_function_conv.scala 1025:26]
  assign sextconv9185_io_enable_bits_taskID = bb_for_body124_io_Out_70_bits_taskID; // @[extracted_function_conv.scala 1025:26]
  assign sextconv9185_io_Out_0_ready = binaryOp_mul9286_io_RightIO_ready; // @[extracted_function_conv.scala 1474:31]
  assign binaryOp_mul9286_clock = clock;
  assign binaryOp_mul9286_reset = reset;
  assign binaryOp_mul9286_io_enable_valid = bb_for_body124_io_Out_71_valid; // @[extracted_function_conv.scala 1028:30]
  assign binaryOp_mul9286_io_enable_bits_taskID = bb_for_body124_io_Out_71_bits_taskID; // @[extracted_function_conv.scala 1028:30]
  assign binaryOp_mul9286_io_enable_bits_control = bb_for_body124_io_Out_71_bits_control; // @[extracted_function_conv.scala 1028:30]
  assign binaryOp_mul9286_io_Out_0_ready = binaryOp_add9387_io_LeftIO_ready; // @[extracted_function_conv.scala 1476:30]
  assign binaryOp_mul9286_io_LeftIO_valid = ld_81_io_Out_0_valid; // @[extracted_function_conv.scala 1462:30]
  assign binaryOp_mul9286_io_LeftIO_bits_data = ld_81_io_Out_0_bits_data; // @[extracted_function_conv.scala 1462:30]
  assign binaryOp_mul9286_io_RightIO_valid = sextconv9185_io_Out_0_valid; // @[extracted_function_conv.scala 1474:31]
  assign binaryOp_mul9286_io_RightIO_bits_data = sextconv9185_io_Out_0_bits_data; // @[extracted_function_conv.scala 1474:31]
  assign binaryOp_add9387_clock = clock;
  assign binaryOp_add9387_reset = reset;
  assign binaryOp_add9387_io_enable_valid = bb_for_body124_io_Out_72_valid; // @[extracted_function_conv.scala 1031:30]
  assign binaryOp_add9387_io_enable_bits_taskID = bb_for_body124_io_Out_72_bits_taskID; // @[extracted_function_conv.scala 1031:30]
  assign binaryOp_add9387_io_enable_bits_control = bb_for_body124_io_Out_72_bits_control; // @[extracted_function_conv.scala 1031:30]
  assign binaryOp_add9387_io_Out_0_ready = st_88_io_inData_ready; // @[extracted_function_conv.scala 1478:19]
  assign binaryOp_add9387_io_Out_1_ready = binaryOp_add10595_io_RightIO_ready; // @[extracted_function_conv.scala 1480:32]
  assign binaryOp_add9387_io_LeftIO_valid = binaryOp_mul9286_io_Out_0_valid; // @[extracted_function_conv.scala 1476:30]
  assign binaryOp_add9387_io_LeftIO_bits_data = binaryOp_mul9286_io_Out_0_bits_data; // @[extracted_function_conv.scala 1476:30]
  assign binaryOp_add9387_io_RightIO_valid = binaryOp_add8279_io_Out_1_valid; // @[extracted_function_conv.scala 1460:31]
  assign binaryOp_add9387_io_RightIO_bits_data = binaryOp_add8279_io_Out_1_bits_data; // @[extracted_function_conv.scala 1460:31]
  assign st_88_clock = clock;
  assign st_88_reset = reset;
  assign st_88_io_enable_valid = bb_for_body124_io_Out_73_valid; // @[extracted_function_conv.scala 1034:19]
  assign st_88_io_enable_bits_taskID = bb_for_body124_io_Out_73_bits_taskID; // @[extracted_function_conv.scala 1034:19]
  assign st_88_io_enable_bits_control = bb_for_body124_io_Out_73_bits_control; // @[extracted_function_conv.scala 1034:19]
  assign st_88_io_GepAddr_valid = Gep_arrayidx28_io_Out_7_valid; // @[extracted_function_conv.scala 1342:20]
  assign st_88_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_7_bits_taskID; // @[extracted_function_conv.scala 1342:20]
  assign st_88_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_7_bits_data; // @[extracted_function_conv.scala 1342:20]
  assign st_88_io_inData_valid = binaryOp_add9387_io_Out_0_valid; // @[extracted_function_conv.scala 1478:19]
  assign st_88_io_inData_bits_taskID = binaryOp_add9387_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1478:19]
  assign st_88_io_inData_bits_data = binaryOp_add9387_io_Out_0_bits_data; // @[extracted_function_conv.scala 1478:19]
  assign st_88_io_memReq_ready = MemCtrl_io_WriteIn_6_ready; // @[extracted_function_conv.scala 1200:25]
  assign st_88_io_memResp_valid = MemCtrl_io_WriteOut_6_valid; // @[extracted_function_conv.scala 1202:20]
  assign ld_89_clock = clock;
  assign ld_89_reset = reset;
  assign ld_89_io_enable_valid = bb_for_body124_io_Out_74_valid; // @[extracted_function_conv.scala 1037:19]
  assign ld_89_io_enable_bits_taskID = bb_for_body124_io_Out_74_bits_taskID; // @[extracted_function_conv.scala 1037:19]
  assign ld_89_io_enable_bits_control = bb_for_body124_io_Out_74_bits_control; // @[extracted_function_conv.scala 1037:19]
  assign ld_89_io_Out_0_ready = binaryOp_mul10494_io_LeftIO_ready; // @[extracted_function_conv.scala 1482:31]
  assign ld_89_io_GepAddr_valid = Loop_0_io_OutLiveIn_field9_0_valid; // @[extracted_function_conv.scala 640:20]
  assign ld_89_io_GepAddr_bits_predicate = Loop_0_io_OutLiveIn_field9_0_bits_predicate; // @[extracted_function_conv.scala 640:20]
  assign ld_89_io_GepAddr_bits_taskID = Loop_0_io_OutLiveIn_field9_0_bits_taskID; // @[extracted_function_conv.scala 640:20]
  assign ld_89_io_GepAddr_bits_data = Loop_0_io_OutLiveIn_field9_0_bits_data; // @[extracted_function_conv.scala 640:20]
  assign ld_89_io_memReq_ready = MemCtrl_io_ReadIn_15_ready; // @[extracted_function_conv.scala 1204:25]
  assign ld_89_io_memResp_valid = MemCtrl_io_ReadOut_15_valid; // @[extracted_function_conv.scala 1206:20]
  assign ld_89_io_memResp_data = MemCtrl_io_ReadOut_15_data; // @[extracted_function_conv.scala 1206:20]
  assign binaryOp_add10090_clock = clock;
  assign binaryOp_add10090_reset = reset;
  assign binaryOp_add10090_io_enable_valid = bb_for_body124_io_Out_75_valid; // @[extracted_function_conv.scala 1040:31]
  assign binaryOp_add10090_io_enable_bits_taskID = bb_for_body124_io_Out_75_bits_taskID; // @[extracted_function_conv.scala 1040:31]
  assign binaryOp_add10090_io_enable_bits_control = bb_for_body124_io_Out_75_bits_control; // @[extracted_function_conv.scala 1040:31]
  assign binaryOp_add10090_io_Out_0_ready = Gep_arrayidx10191_io_idx_0_ready; // @[extracted_function_conv.scala 1484:31]
  assign binaryOp_add10090_io_LeftIO_valid = binaryOp_add8882_io_Out_1_valid; // @[extracted_function_conv.scala 1466:31]
  assign binaryOp_add10090_io_LeftIO_bits_data = binaryOp_add8882_io_Out_1_bits_data; // @[extracted_function_conv.scala 1466:31]
  assign binaryOp_add10090_io_RightIO_valid = const22_io_Out_valid; // @[extracted_function_conv.scala 1284:32]
  assign Gep_arrayidx10191_clock = clock;
  assign Gep_arrayidx10191_reset = reset;
  assign Gep_arrayidx10191_io_enable_valid = bb_for_body124_io_Out_76_valid; // @[extracted_function_conv.scala 1043:31]
  assign Gep_arrayidx10191_io_enable_bits_taskID = bb_for_body124_io_Out_76_bits_taskID; // @[extracted_function_conv.scala 1043:31]
  assign Gep_arrayidx10191_io_enable_bits_control = bb_for_body124_io_Out_76_bits_control; // @[extracted_function_conv.scala 1043:31]
  assign Gep_arrayidx10191_io_Out_0_ready = ld_92_io_GepAddr_ready; // @[extracted_function_conv.scala 1486:20]
  assign Gep_arrayidx10191_io_baseAddress_valid = Loop_0_io_OutLiveIn_field10_7_valid; // @[extracted_function_conv.scala 656:36]
  assign Gep_arrayidx10191_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field10_7_bits_taskID; // @[extracted_function_conv.scala 656:36]
  assign Gep_arrayidx10191_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field10_7_bits_data; // @[extracted_function_conv.scala 656:36]
  assign Gep_arrayidx10191_io_idx_0_valid = binaryOp_add10090_io_Out_0_valid; // @[extracted_function_conv.scala 1484:31]
  assign Gep_arrayidx10191_io_idx_0_bits_data = binaryOp_add10090_io_Out_0_bits_data; // @[extracted_function_conv.scala 1484:31]
  assign ld_92_clock = clock;
  assign ld_92_reset = reset;
  assign ld_92_io_enable_valid = bb_for_body124_io_Out_77_valid; // @[extracted_function_conv.scala 1046:19]
  assign ld_92_io_enable_bits_taskID = bb_for_body124_io_Out_77_bits_taskID; // @[extracted_function_conv.scala 1046:19]
  assign ld_92_io_enable_bits_control = bb_for_body124_io_Out_77_bits_control; // @[extracted_function_conv.scala 1046:19]
  assign ld_92_io_Out_0_ready = sextconv10393_io_Input_ready; // @[extracted_function_conv.scala 1488:26]
  assign ld_92_io_GepAddr_valid = Gep_arrayidx10191_io_Out_0_valid; // @[extracted_function_conv.scala 1486:20]
  assign ld_92_io_GepAddr_bits_predicate = Gep_arrayidx10191_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1486:20]
  assign ld_92_io_GepAddr_bits_taskID = Gep_arrayidx10191_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1486:20]
  assign ld_92_io_GepAddr_bits_data = Gep_arrayidx10191_io_Out_0_bits_data; // @[extracted_function_conv.scala 1486:20]
  assign ld_92_io_memReq_ready = MemCtrl_io_ReadIn_16_ready; // @[extracted_function_conv.scala 1208:25]
  assign ld_92_io_memResp_valid = MemCtrl_io_ReadOut_16_valid; // @[extracted_function_conv.scala 1210:20]
  assign ld_92_io_memResp_data = MemCtrl_io_ReadOut_16_data; // @[extracted_function_conv.scala 1210:20]
  assign sextconv10393_clock = clock;
  assign sextconv10393_reset = reset;
  assign sextconv10393_io_Input_valid = ld_92_io_Out_0_valid; // @[extracted_function_conv.scala 1488:26]
  assign sextconv10393_io_Input_bits_data = ld_92_io_Out_0_bits_data; // @[extracted_function_conv.scala 1488:26]
  assign sextconv10393_io_enable_valid = bb_for_body124_io_Out_78_valid; // @[extracted_function_conv.scala 1049:27]
  assign sextconv10393_io_enable_bits_taskID = bb_for_body124_io_Out_78_bits_taskID; // @[extracted_function_conv.scala 1049:27]
  assign sextconv10393_io_Out_0_ready = binaryOp_mul10494_io_RightIO_ready; // @[extracted_function_conv.scala 1490:32]
  assign binaryOp_mul10494_clock = clock;
  assign binaryOp_mul10494_reset = reset;
  assign binaryOp_mul10494_io_enable_valid = bb_for_body124_io_Out_79_valid; // @[extracted_function_conv.scala 1052:31]
  assign binaryOp_mul10494_io_enable_bits_taskID = bb_for_body124_io_Out_79_bits_taskID; // @[extracted_function_conv.scala 1052:31]
  assign binaryOp_mul10494_io_enable_bits_control = bb_for_body124_io_Out_79_bits_control; // @[extracted_function_conv.scala 1052:31]
  assign binaryOp_mul10494_io_Out_0_ready = binaryOp_add10595_io_LeftIO_ready; // @[extracted_function_conv.scala 1492:31]
  assign binaryOp_mul10494_io_LeftIO_valid = ld_89_io_Out_0_valid; // @[extracted_function_conv.scala 1482:31]
  assign binaryOp_mul10494_io_LeftIO_bits_data = ld_89_io_Out_0_bits_data; // @[extracted_function_conv.scala 1482:31]
  assign binaryOp_mul10494_io_RightIO_valid = sextconv10393_io_Out_0_valid; // @[extracted_function_conv.scala 1490:32]
  assign binaryOp_mul10494_io_RightIO_bits_data = sextconv10393_io_Out_0_bits_data; // @[extracted_function_conv.scala 1490:32]
  assign binaryOp_add10595_clock = clock;
  assign binaryOp_add10595_reset = reset;
  assign binaryOp_add10595_io_enable_valid = bb_for_body124_io_Out_80_valid; // @[extracted_function_conv.scala 1055:31]
  assign binaryOp_add10595_io_enable_bits_taskID = bb_for_body124_io_Out_80_bits_taskID; // @[extracted_function_conv.scala 1055:31]
  assign binaryOp_add10595_io_enable_bits_control = bb_for_body124_io_Out_80_bits_control; // @[extracted_function_conv.scala 1055:31]
  assign binaryOp_add10595_io_Out_0_ready = st_96_io_inData_ready; // @[extracted_function_conv.scala 1494:19]
  assign binaryOp_add10595_io_Out_1_ready = binaryOp_add117103_io_RightIO_ready; // @[extracted_function_conv.scala 1496:33]
  assign binaryOp_add10595_io_LeftIO_valid = binaryOp_mul10494_io_Out_0_valid; // @[extracted_function_conv.scala 1492:31]
  assign binaryOp_add10595_io_LeftIO_bits_data = binaryOp_mul10494_io_Out_0_bits_data; // @[extracted_function_conv.scala 1492:31]
  assign binaryOp_add10595_io_RightIO_valid = binaryOp_add9387_io_Out_1_valid; // @[extracted_function_conv.scala 1480:32]
  assign binaryOp_add10595_io_RightIO_bits_data = binaryOp_add9387_io_Out_1_bits_data; // @[extracted_function_conv.scala 1480:32]
  assign st_96_clock = clock;
  assign st_96_reset = reset;
  assign st_96_io_enable_valid = bb_for_body124_io_Out_81_valid; // @[extracted_function_conv.scala 1058:19]
  assign st_96_io_enable_bits_taskID = bb_for_body124_io_Out_81_bits_taskID; // @[extracted_function_conv.scala 1058:19]
  assign st_96_io_enable_bits_control = bb_for_body124_io_Out_81_bits_control; // @[extracted_function_conv.scala 1058:19]
  assign st_96_io_GepAddr_valid = Gep_arrayidx28_io_Out_8_valid; // @[extracted_function_conv.scala 1344:20]
  assign st_96_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_8_bits_taskID; // @[extracted_function_conv.scala 1344:20]
  assign st_96_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_8_bits_data; // @[extracted_function_conv.scala 1344:20]
  assign st_96_io_inData_valid = binaryOp_add10595_io_Out_0_valid; // @[extracted_function_conv.scala 1494:19]
  assign st_96_io_inData_bits_taskID = binaryOp_add10595_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1494:19]
  assign st_96_io_inData_bits_data = binaryOp_add10595_io_Out_0_bits_data; // @[extracted_function_conv.scala 1494:19]
  assign st_96_io_memReq_ready = MemCtrl_io_WriteIn_7_ready; // @[extracted_function_conv.scala 1212:25]
  assign st_96_io_memResp_valid = MemCtrl_io_WriteOut_7_valid; // @[extracted_function_conv.scala 1214:20]
  assign ld_97_clock = clock;
  assign ld_97_reset = reset;
  assign ld_97_io_enable_valid = bb_for_body124_io_Out_82_valid; // @[extracted_function_conv.scala 1061:19]
  assign ld_97_io_enable_bits_taskID = bb_for_body124_io_Out_82_bits_taskID; // @[extracted_function_conv.scala 1061:19]
  assign ld_97_io_enable_bits_control = bb_for_body124_io_Out_82_bits_control; // @[extracted_function_conv.scala 1061:19]
  assign ld_97_io_Out_0_ready = binaryOp_mul116102_io_LeftIO_ready; // @[extracted_function_conv.scala 1498:32]
  assign ld_97_io_GepAddr_valid = Loop_0_io_OutLiveIn_field4_0_valid; // @[extracted_function_conv.scala 630:20]
  assign ld_97_io_GepAddr_bits_predicate = Loop_0_io_OutLiveIn_field4_0_bits_predicate; // @[extracted_function_conv.scala 630:20]
  assign ld_97_io_GepAddr_bits_taskID = Loop_0_io_OutLiveIn_field4_0_bits_taskID; // @[extracted_function_conv.scala 630:20]
  assign ld_97_io_GepAddr_bits_data = Loop_0_io_OutLiveIn_field4_0_bits_data; // @[extracted_function_conv.scala 630:20]
  assign ld_97_io_memReq_ready = MemCtrl_io_ReadIn_17_ready; // @[extracted_function_conv.scala 1216:25]
  assign ld_97_io_memResp_valid = MemCtrl_io_ReadOut_17_valid; // @[extracted_function_conv.scala 1218:20]
  assign ld_97_io_memResp_data = MemCtrl_io_ReadOut_17_data; // @[extracted_function_conv.scala 1218:20]
  assign binaryOp_add11298_clock = clock;
  assign binaryOp_add11298_reset = reset;
  assign binaryOp_add11298_io_enable_valid = bb_for_body124_io_Out_83_valid; // @[extracted_function_conv.scala 1064:31]
  assign binaryOp_add11298_io_enable_bits_taskID = bb_for_body124_io_Out_83_bits_taskID; // @[extracted_function_conv.scala 1064:31]
  assign binaryOp_add11298_io_enable_bits_control = bb_for_body124_io_Out_83_bits_control; // @[extracted_function_conv.scala 1064:31]
  assign binaryOp_add11298_io_Out_0_ready = Gep_arrayidx11399_io_idx_0_ready; // @[extracted_function_conv.scala 1500:31]
  assign binaryOp_add11298_io_LeftIO_valid = binaryOp_add8882_io_Out_2_valid; // @[extracted_function_conv.scala 1468:31]
  assign binaryOp_add11298_io_LeftIO_bits_data = binaryOp_add8882_io_Out_2_bits_data; // @[extracted_function_conv.scala 1468:31]
  assign binaryOp_add11298_io_RightIO_valid = const23_io_Out_valid; // @[extracted_function_conv.scala 1286:32]
  assign Gep_arrayidx11399_clock = clock;
  assign Gep_arrayidx11399_reset = reset;
  assign Gep_arrayidx11399_io_enable_valid = bb_for_body124_io_Out_84_valid; // @[extracted_function_conv.scala 1067:31]
  assign Gep_arrayidx11399_io_enable_bits_taskID = bb_for_body124_io_Out_84_bits_taskID; // @[extracted_function_conv.scala 1067:31]
  assign Gep_arrayidx11399_io_enable_bits_control = bb_for_body124_io_Out_84_bits_control; // @[extracted_function_conv.scala 1067:31]
  assign Gep_arrayidx11399_io_Out_0_ready = ld_100_io_GepAddr_ready; // @[extracted_function_conv.scala 1502:21]
  assign Gep_arrayidx11399_io_baseAddress_valid = Loop_0_io_OutLiveIn_field10_8_valid; // @[extracted_function_conv.scala 658:36]
  assign Gep_arrayidx11399_io_baseAddress_bits_taskID = Loop_0_io_OutLiveIn_field10_8_bits_taskID; // @[extracted_function_conv.scala 658:36]
  assign Gep_arrayidx11399_io_baseAddress_bits_data = Loop_0_io_OutLiveIn_field10_8_bits_data; // @[extracted_function_conv.scala 658:36]
  assign Gep_arrayidx11399_io_idx_0_valid = binaryOp_add11298_io_Out_0_valid; // @[extracted_function_conv.scala 1500:31]
  assign Gep_arrayidx11399_io_idx_0_bits_data = binaryOp_add11298_io_Out_0_bits_data; // @[extracted_function_conv.scala 1500:31]
  assign ld_100_clock = clock;
  assign ld_100_reset = reset;
  assign ld_100_io_enable_valid = bb_for_body124_io_Out_85_valid; // @[extracted_function_conv.scala 1070:20]
  assign ld_100_io_enable_bits_taskID = bb_for_body124_io_Out_85_bits_taskID; // @[extracted_function_conv.scala 1070:20]
  assign ld_100_io_enable_bits_control = bb_for_body124_io_Out_85_bits_control; // @[extracted_function_conv.scala 1070:20]
  assign ld_100_io_Out_0_ready = sextconv115101_io_Input_ready; // @[extracted_function_conv.scala 1504:27]
  assign ld_100_io_GepAddr_valid = Gep_arrayidx11399_io_Out_0_valid; // @[extracted_function_conv.scala 1502:21]
  assign ld_100_io_GepAddr_bits_predicate = Gep_arrayidx11399_io_Out_0_bits_predicate; // @[extracted_function_conv.scala 1502:21]
  assign ld_100_io_GepAddr_bits_taskID = Gep_arrayidx11399_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1502:21]
  assign ld_100_io_GepAddr_bits_data = Gep_arrayidx11399_io_Out_0_bits_data; // @[extracted_function_conv.scala 1502:21]
  assign ld_100_io_memReq_ready = MemCtrl_io_ReadIn_18_ready; // @[extracted_function_conv.scala 1220:25]
  assign ld_100_io_memResp_valid = MemCtrl_io_ReadOut_18_valid; // @[extracted_function_conv.scala 1222:21]
  assign ld_100_io_memResp_data = MemCtrl_io_ReadOut_18_data; // @[extracted_function_conv.scala 1222:21]
  assign sextconv115101_clock = clock;
  assign sextconv115101_reset = reset;
  assign sextconv115101_io_Input_valid = ld_100_io_Out_0_valid; // @[extracted_function_conv.scala 1504:27]
  assign sextconv115101_io_Input_bits_data = ld_100_io_Out_0_bits_data; // @[extracted_function_conv.scala 1504:27]
  assign sextconv115101_io_enable_valid = bb_for_body124_io_Out_86_valid; // @[extracted_function_conv.scala 1073:28]
  assign sextconv115101_io_enable_bits_taskID = bb_for_body124_io_Out_86_bits_taskID; // @[extracted_function_conv.scala 1073:28]
  assign sextconv115101_io_Out_0_ready = binaryOp_mul116102_io_RightIO_ready; // @[extracted_function_conv.scala 1506:33]
  assign binaryOp_mul116102_clock = clock;
  assign binaryOp_mul116102_reset = reset;
  assign binaryOp_mul116102_io_enable_valid = bb_for_body124_io_Out_87_valid; // @[extracted_function_conv.scala 1076:32]
  assign binaryOp_mul116102_io_enable_bits_taskID = bb_for_body124_io_Out_87_bits_taskID; // @[extracted_function_conv.scala 1076:32]
  assign binaryOp_mul116102_io_enable_bits_control = bb_for_body124_io_Out_87_bits_control; // @[extracted_function_conv.scala 1076:32]
  assign binaryOp_mul116102_io_Out_0_ready = binaryOp_add117103_io_LeftIO_ready; // @[extracted_function_conv.scala 1508:32]
  assign binaryOp_mul116102_io_LeftIO_valid = ld_97_io_Out_0_valid; // @[extracted_function_conv.scala 1498:32]
  assign binaryOp_mul116102_io_LeftIO_bits_data = ld_97_io_Out_0_bits_data; // @[extracted_function_conv.scala 1498:32]
  assign binaryOp_mul116102_io_RightIO_valid = sextconv115101_io_Out_0_valid; // @[extracted_function_conv.scala 1506:33]
  assign binaryOp_mul116102_io_RightIO_bits_data = sextconv115101_io_Out_0_bits_data; // @[extracted_function_conv.scala 1506:33]
  assign binaryOp_add117103_clock = clock;
  assign binaryOp_add117103_reset = reset;
  assign binaryOp_add117103_io_enable_valid = bb_for_body124_io_Out_88_valid; // @[extracted_function_conv.scala 1079:32]
  assign binaryOp_add117103_io_enable_bits_taskID = bb_for_body124_io_Out_88_bits_taskID; // @[extracted_function_conv.scala 1079:32]
  assign binaryOp_add117103_io_enable_bits_control = bb_for_body124_io_Out_88_bits_control; // @[extracted_function_conv.scala 1079:32]
  assign binaryOp_add117103_io_Out_0_ready = st_104_io_inData_ready; // @[extracted_function_conv.scala 1510:20]
  assign binaryOp_add117103_io_LeftIO_valid = binaryOp_mul116102_io_Out_0_valid; // @[extracted_function_conv.scala 1508:32]
  assign binaryOp_add117103_io_LeftIO_bits_data = binaryOp_mul116102_io_Out_0_bits_data; // @[extracted_function_conv.scala 1508:32]
  assign binaryOp_add117103_io_RightIO_valid = binaryOp_add10595_io_Out_1_valid; // @[extracted_function_conv.scala 1496:33]
  assign binaryOp_add117103_io_RightIO_bits_data = binaryOp_add10595_io_Out_1_bits_data; // @[extracted_function_conv.scala 1496:33]
  assign st_104_clock = clock;
  assign st_104_reset = reset;
  assign st_104_io_enable_valid = bb_for_body124_io_Out_89_valid; // @[extracted_function_conv.scala 1082:20]
  assign st_104_io_enable_bits_taskID = bb_for_body124_io_Out_89_bits_taskID; // @[extracted_function_conv.scala 1082:20]
  assign st_104_io_enable_bits_control = bb_for_body124_io_Out_89_bits_control; // @[extracted_function_conv.scala 1082:20]
  assign st_104_io_GepAddr_valid = Gep_arrayidx28_io_Out_9_valid; // @[extracted_function_conv.scala 1346:21]
  assign st_104_io_GepAddr_bits_taskID = Gep_arrayidx28_io_Out_9_bits_taskID; // @[extracted_function_conv.scala 1346:21]
  assign st_104_io_GepAddr_bits_data = Gep_arrayidx28_io_Out_9_bits_data; // @[extracted_function_conv.scala 1346:21]
  assign st_104_io_inData_valid = binaryOp_add117103_io_Out_0_valid; // @[extracted_function_conv.scala 1510:20]
  assign st_104_io_inData_bits_taskID = binaryOp_add117103_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1510:20]
  assign st_104_io_inData_bits_data = binaryOp_add117103_io_Out_0_bits_data; // @[extracted_function_conv.scala 1510:20]
  assign st_104_io_memReq_ready = MemCtrl_io_WriteIn_8_ready; // @[extracted_function_conv.scala 1224:25]
  assign st_104_io_memResp_valid = MemCtrl_io_WriteOut_8_valid; // @[extracted_function_conv.scala 1226:21]
  assign binaryOp_inc105_clock = clock;
  assign binaryOp_inc105_reset = reset;
  assign binaryOp_inc105_io_enable_valid = bb_for_body124_io_Out_90_valid; // @[extracted_function_conv.scala 1085:29]
  assign binaryOp_inc105_io_enable_bits_taskID = bb_for_body124_io_Out_90_bits_taskID; // @[extracted_function_conv.scala 1085:29]
  assign binaryOp_inc105_io_enable_bits_control = bb_for_body124_io_Out_90_bits_control; // @[extracted_function_conv.scala 1085:29]
  assign binaryOp_inc105_io_Out_0_ready = Loop_0_io_CarryDepenIn_0_ready; // @[extracted_function_conv.scala 698:29]
  assign binaryOp_inc105_io_Out_1_ready = icmp_exitcond106_io_LeftIO_ready; // @[extracted_function_conv.scala 1512:30]
  assign binaryOp_inc105_io_LeftIO_valid = phi_conv_s1_x_031226_io_Out_3_valid; // @[extracted_function_conv.scala 1324:29]
  assign binaryOp_inc105_io_LeftIO_bits_data = phi_conv_s1_x_031226_io_Out_3_bits_data; // @[extracted_function_conv.scala 1324:29]
  assign binaryOp_inc105_io_RightIO_valid = const24_io_Out_valid; // @[extracted_function_conv.scala 1288:30]
  assign icmp_exitcond106_clock = clock;
  assign icmp_exitcond106_reset = reset;
  assign icmp_exitcond106_io_enable_valid = bb_for_body124_io_Out_91_valid; // @[extracted_function_conv.scala 1088:30]
  assign icmp_exitcond106_io_enable_bits_taskID = bb_for_body124_io_Out_91_bits_taskID; // @[extracted_function_conv.scala 1088:30]
  assign icmp_exitcond106_io_enable_bits_control = bb_for_body124_io_Out_91_bits_control; // @[extracted_function_conv.scala 1088:30]
  assign icmp_exitcond106_io_Out_0_ready = br_107_io_CmpIO_ready; // @[extracted_function_conv.scala 1514:19]
  assign icmp_exitcond106_io_LeftIO_valid = binaryOp_inc105_io_Out_1_valid; // @[extracted_function_conv.scala 1512:30]
  assign icmp_exitcond106_io_LeftIO_bits_data = binaryOp_inc105_io_Out_1_bits_data; // @[extracted_function_conv.scala 1512:30]
  assign icmp_exitcond106_io_RightIO_valid = const25_io_Out_valid; // @[extracted_function_conv.scala 1290:31]
  assign br_107_clock = clock;
  assign br_107_reset = reset;
  assign br_107_io_enable_valid = bb_for_body124_io_Out_92_valid; // @[extracted_function_conv.scala 1091:20]
  assign br_107_io_enable_bits_taskID = bb_for_body124_io_Out_92_bits_taskID; // @[extracted_function_conv.scala 1091:20]
  assign br_107_io_enable_bits_control = bb_for_body124_io_Out_92_bits_control; // @[extracted_function_conv.scala 1091:20]
  assign br_107_io_CmpIO_valid = icmp_exitcond106_io_Out_0_valid; // @[extracted_function_conv.scala 1514:19]
  assign br_107_io_CmpIO_bits_taskID = icmp_exitcond106_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 1514:19]
  assign br_107_io_CmpIO_bits_data = icmp_exitcond106_io_Out_0_bits_data; // @[extracted_function_conv.scala 1514:19]
  assign br_107_io_TrueOutput_0_ready = Loop_0_io_loopFinish_0_ready; // @[extracted_function_conv.scala 538:27]
  assign br_107_io_FalseOutput_0_ready = Loop_0_io_loopBack_0_ready; // @[extracted_function_conv.scala 536:25]
  assign const0_clock = clock;
  assign const0_reset = reset;
  assign const0_io_enable_valid = bb_entry0_io_Out_0_valid; // @[extracted_function_conv.scala 718:20]
  assign const0_io_enable_bits_taskID = bb_entry0_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 718:20]
  assign const0_io_Out_ready = Gep_arrayidx252_io_idx_0_ready; // @[extracted_function_conv.scala 1240:29]
  assign const1_clock = clock;
  assign const1_reset = reset;
  assign const1_io_enable_valid = bb_entry0_io_Out_1_valid; // @[extracted_function_conv.scala 720:20]
  assign const1_io_enable_bits_taskID = bb_entry0_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 720:20]
  assign const1_io_Out_ready = Gep_arrayidx383_io_idx_0_ready; // @[extracted_function_conv.scala 1242:29]
  assign const2_clock = clock;
  assign const2_reset = reset;
  assign const2_io_enable_valid = bb_entry0_io_Out_2_valid; // @[extracted_function_conv.scala 722:20]
  assign const2_io_enable_bits_taskID = bb_entry0_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 722:20]
  assign const2_io_Out_ready = Gep_arrayidx514_io_idx_0_ready; // @[extracted_function_conv.scala 1244:29]
  assign const3_clock = clock;
  assign const3_reset = reset;
  assign const3_io_enable_valid = bb_entry0_io_Out_3_valid; // @[extracted_function_conv.scala 724:20]
  assign const3_io_enable_bits_taskID = bb_entry0_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 724:20]
  assign const3_io_Out_ready = Gep_arrayidx625_io_idx_0_ready; // @[extracted_function_conv.scala 1246:29]
  assign const4_clock = clock;
  assign const4_reset = reset;
  assign const4_io_enable_valid = bb_entry0_io_Out_4_valid; // @[extracted_function_conv.scala 726:20]
  assign const4_io_enable_bits_taskID = bb_entry0_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 726:20]
  assign const4_io_Out_ready = Gep_arrayidx746_io_idx_0_ready; // @[extracted_function_conv.scala 1248:29]
  assign const5_clock = clock;
  assign const5_reset = reset;
  assign const5_io_enable_valid = bb_entry0_io_Out_5_valid; // @[extracted_function_conv.scala 728:20]
  assign const5_io_enable_bits_taskID = bb_entry0_io_Out_5_bits_taskID; // @[extracted_function_conv.scala 728:20]
  assign const5_io_Out_ready = Gep_arrayidx867_io_idx_0_ready; // @[extracted_function_conv.scala 1250:29]
  assign const6_clock = clock;
  assign const6_reset = reset;
  assign const6_io_enable_valid = bb_entry0_io_Out_6_valid; // @[extracted_function_conv.scala 730:20]
  assign const6_io_enable_bits_taskID = bb_entry0_io_Out_6_bits_taskID; // @[extracted_function_conv.scala 730:20]
  assign const6_io_Out_ready = Gep_arrayidx978_io_idx_0_ready; // @[extracted_function_conv.scala 1252:29]
  assign const7_clock = clock;
  assign const7_reset = reset;
  assign const7_io_enable_valid = bb_entry0_io_Out_7_valid; // @[extracted_function_conv.scala 732:20]
  assign const7_io_enable_bits_taskID = bb_entry0_io_Out_7_bits_taskID; // @[extracted_function_conv.scala 732:20]
  assign const7_io_Out_ready = Gep_arrayidx1099_io_idx_0_ready; // @[extracted_function_conv.scala 1254:30]
  assign const8_clock = clock;
  assign const8_reset = reset;
  assign const8_io_enable_valid = bb_for_body2_io_Out_0_valid; // @[extracted_function_conv.scala 770:20]
  assign const8_io_enable_bits_taskID = bb_for_body2_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 770:20]
  assign const8_io_Out_ready = phi_conv_s1_y_031312_io_InData_0_ready; // @[extracted_function_conv.scala 1256:37]
  assign const9_clock = clock;
  assign const9_reset = reset;
  assign const9_io_enable_valid = bb_for_body2_io_Out_1_valid; // @[extracted_function_conv.scala 772:20]
  assign const9_io_enable_bits_taskID = bb_for_body2_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 772:20]
  assign const9_io_Out_ready = binaryOp_mul113_io_RightIO_ready; // @[extracted_function_conv.scala 1258:30]
  assign const10_clock = clock;
  assign const10_reset = reset;
  assign const10_io_enable_valid = bb_for_body2_io_Out_2_valid; // @[extracted_function_conv.scala 774:21]
  assign const10_io_enable_bits_taskID = bb_for_body2_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 774:21]
  assign const10_io_Out_ready = binaryOp_add214_io_RightIO_ready; // @[extracted_function_conv.scala 1260:30]
  assign const11_clock = clock;
  assign const11_reset = reset;
  assign const11_io_enable_valid = bb_for_body2_io_Out_3_valid; // @[extracted_function_conv.scala 776:21]
  assign const11_io_enable_bits_taskID = bb_for_body2_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 776:21]
  assign const11_io_Out_ready = binaryOp_add417_io_RightIO_ready; // @[extracted_function_conv.scala 1262:30]
  assign const12_clock = clock;
  assign const12_reset = reset;
  assign const12_io_enable_valid = bb_for_body2_io_Out_4_valid; // @[extracted_function_conv.scala 778:21]
  assign const12_io_enable_bits_taskID = bb_for_body2_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 778:21]
  assign const12_io_Out_ready = binaryOp_mul821_io_RightIO_ready; // @[extracted_function_conv.scala 1264:30]
  assign const13_clock = clock;
  assign const13_reset = reset;
  assign const13_io_enable_valid = bb_for_cond_cleanup113_io_Out_0_valid; // @[extracted_function_conv.scala 813:21]
  assign const13_io_enable_bits_taskID = bb_for_cond_cleanup113_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 813:21]
  assign const13_io_Out_ready = binaryOp_inc12023_io_RightIO_ready; // @[extracted_function_conv.scala 1266:32]
  assign const14_clock = clock;
  assign const14_reset = reset;
  assign const14_io_enable_valid = bb_for_cond_cleanup113_io_Out_1_valid; // @[extracted_function_conv.scala 815:21]
  assign const14_io_enable_bits_taskID = bb_for_cond_cleanup113_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 815:21]
  assign const14_io_Out_ready = icmp_exitcond31424_io_RightIO_ready; // @[extracted_function_conv.scala 1268:33]
  assign const15_clock = clock;
  assign const15_reset = reset;
  assign const15_io_enable_valid = bb_for_body124_io_Out_0_valid; // @[extracted_function_conv.scala 826:21]
  assign const15_io_enable_bits_taskID = bb_for_body124_io_Out_0_bits_taskID; // @[extracted_function_conv.scala 826:21]
  assign const15_io_Out_ready = phi_conv_s1_x_031226_io_InData_0_ready; // @[extracted_function_conv.scala 1270:37]
  assign const16_clock = clock;
  assign const16_reset = reset;
  assign const16_io_enable_valid = bb_for_body124_io_Out_1_valid; // @[extracted_function_conv.scala 828:21]
  assign const16_io_enable_bits_taskID = bb_for_body124_io_Out_1_bits_taskID; // @[extracted_function_conv.scala 828:21]
  assign const16_io_Out_ready = binaryOp_mul1632_io_RightIO_ready; // @[extracted_function_conv.scala 1272:31]
  assign const17_clock = clock;
  assign const17_reset = reset;
  assign const17_io_enable_valid = bb_for_body124_io_Out_2_valid; // @[extracted_function_conv.scala 830:21]
  assign const17_io_enable_bits_taskID = bb_for_body124_io_Out_2_bits_taskID; // @[extracted_function_conv.scala 830:21]
  assign const17_io_Out_ready = binaryOp_add2941_io_RightIO_ready; // @[extracted_function_conv.scala 1274:31]
  assign const18_clock = clock;
  assign const18_reset = reset;
  assign const18_io_enable_valid = bb_for_body124_io_Out_3_valid; // @[extracted_function_conv.scala 832:21]
  assign const18_io_enable_bits_taskID = bb_for_body124_io_Out_3_bits_taskID; // @[extracted_function_conv.scala 832:21]
  assign const18_io_Out_ready = binaryOp_add4249_io_RightIO_ready; // @[extracted_function_conv.scala 1276:31]
  assign const19_clock = clock;
  assign const19_reset = reset;
  assign const19_io_enable_valid = bb_for_body124_io_Out_4_valid; // @[extracted_function_conv.scala 834:21]
  assign const19_io_enable_bits_taskID = bb_for_body124_io_Out_4_bits_taskID; // @[extracted_function_conv.scala 834:21]
  assign const19_io_Out_ready = binaryOp_mul5257_io_RightIO_ready; // @[extracted_function_conv.scala 1278:31]
  assign const20_clock = clock;
  assign const20_reset = reset;
  assign const20_io_enable_valid = bb_for_body124_io_Out_5_valid; // @[extracted_function_conv.scala 836:21]
  assign const20_io_enable_bits_taskID = bb_for_body124_io_Out_5_bits_taskID; // @[extracted_function_conv.scala 836:21]
  assign const20_io_Out_ready = binaryOp_add6566_io_RightIO_ready; // @[extracted_function_conv.scala 1280:31]
  assign const21_clock = clock;
  assign const21_reset = reset;
  assign const21_io_enable_valid = bb_for_body124_io_Out_6_valid; // @[extracted_function_conv.scala 838:21]
  assign const21_io_enable_bits_taskID = bb_for_body124_io_Out_6_bits_taskID; // @[extracted_function_conv.scala 838:21]
  assign const21_io_Out_ready = binaryOp_add7774_io_RightIO_ready; // @[extracted_function_conv.scala 1282:31]
  assign const22_clock = clock;
  assign const22_reset = reset;
  assign const22_io_enable_valid = bb_for_body124_io_Out_7_valid; // @[extracted_function_conv.scala 840:21]
  assign const22_io_enable_bits_taskID = bb_for_body124_io_Out_7_bits_taskID; // @[extracted_function_conv.scala 840:21]
  assign const22_io_Out_ready = binaryOp_add10090_io_RightIO_ready; // @[extracted_function_conv.scala 1284:32]
  assign const23_clock = clock;
  assign const23_reset = reset;
  assign const23_io_enable_valid = bb_for_body124_io_Out_8_valid; // @[extracted_function_conv.scala 842:21]
  assign const23_io_enable_bits_taskID = bb_for_body124_io_Out_8_bits_taskID; // @[extracted_function_conv.scala 842:21]
  assign const23_io_Out_ready = binaryOp_add11298_io_RightIO_ready; // @[extracted_function_conv.scala 1286:32]
  assign const24_clock = clock;
  assign const24_reset = reset;
  assign const24_io_enable_valid = bb_for_body124_io_Out_9_valid; // @[extracted_function_conv.scala 844:21]
  assign const24_io_enable_bits_taskID = bb_for_body124_io_Out_9_bits_taskID; // @[extracted_function_conv.scala 844:21]
  assign const24_io_Out_ready = binaryOp_inc105_io_RightIO_ready; // @[extracted_function_conv.scala 1288:30]
  assign const25_clock = clock;
  assign const25_reset = reset;
  assign const25_io_enable_valid = bb_for_body124_io_Out_10_valid; // @[extracted_function_conv.scala 846:21]
  assign const25_io_enable_bits_taskID = bb_for_body124_io_Out_10_bits_taskID; // @[extracted_function_conv.scala 846:21]
  assign const25_io_Out_ready = icmp_exitcond106_io_RightIO_ready; // @[extracted_function_conv.scala 1290:31]
endmodule
